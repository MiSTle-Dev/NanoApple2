--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.10.03 (64-bit)
--Part Number: GW5AT-LV60PG484AC1/I0
--Device: GW5AT-60
--Device Version: B
--Created Time: Tue May 27 15:16:48 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_video is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(11 downto 0)
    );
end Gowin_pROM_video;

architecture Behavioral of Gowin_pROM_video is

    signal prom_inst_0_dout_w: std_logic_vector(27 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(27 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(3 downto 0) <= prom_inst_0_DO_o(3 downto 0) ;
    prom_inst_0_dout_w(27 downto 0) <= prom_inst_0_DO_o(31 downto 4) ;
    prom_inst_1_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(7 downto 4) <= prom_inst_1_DO_o(3 downto 0) ;
    prom_inst_1_dout_w(27 downto 0) <= prom_inst_1_DO_o(31 downto 4) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 4,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0C22222C0222E22E0E22E22E0E22222E0C22222C0E22E22E022E22480C2AAA2C",
            INIT_RAM_01 => X"0C22222C0222A6220222AA620E222222022A6A220C2000000C88888C0222E222",
            INIT_RAM_02 => X"026AA222084222220C2222220888888E0C20C22C022AE22E0C2A222C0222E22E",
            INIT_RAM_03 => X"F0000000000248000E00000E000084200E66666E0E24800E0888842202248422",
            INIT_RAM_04 => X"000008880C2A4AA40024806608E8CAC80A44E448000004440808888800000000",
            INIT_RAM_05 => X"00248000080000000000E000048800000088E88008AC8CA80800000808422248",
            INIT_RAM_06 => X"0444800E0C22E2480C200E2E000E24800C20800E0E24802C0C8888C80C26A22C",
            INIT_RAM_07 => X"0808802C04800084000E0E000084248004880800000808000E00C22C0C22C22C",
            INIT_RAM_08 => X"F738F87FD0F6E1FF044A3000FBB5EFFF05B77BD0D9119DFF95EEE97F9100097F",
            INIT_RAM_09 => X"0F73137C00000000B909BFFFFFFFFFF077776537735677775FFFFFFFF7BD0DB7",
            INIT_RAM_0A => X"5A5A5A5AA5A5A5A5F7FF0FF70EEEEEEEFFFF0FFFF770137FF731077F4B33033B",
            INIT_RAM_0B => X"EEEEEEEE0FF33FF0FBB8F8BB0FFFFFF0F7310137FFFFFFFFF0FFF0FFF0EEEE1F",
            INIT_RAM_0C => X"C0C22C000444E4480C2E2C000C222C000C222C000E222E220C2C0C0000000084",
            INIT_RAM_0D => X"0C222C0002222E0002AAA6000C88888C022E2222C20008000C888C0802222E22",
            INIT_RAM_0E => X"06AA2200084222000C22220008444E440E0C2C0002226A0000C22C0022E22E00",
            INIT_RAM_0F => X"00A4A4A0000000AC0E88088E8888888808CC6CC80E480E00C0C2220002484200",
            INIT_RAM_10 => X"F3DDDDD3FDDD1DD1F1DD1DD1F1DDDDD1F3DDDDD3F1DD1DD1FDD1DDB7F3D555D3",
            INIT_RAM_11 => X"F3DDDDD3FDDD59DDFDDD559DF1DDDDDDFDD595DDF3DFFFFFF3777773FDDD1DDD",
            INIT_RAM_12 => X"FD955DDDF7BDDDDDF3DDDDDDF7777771F3DF3DD3FDD51DD1F3D5DDD3FDDD1DD1",
            INIT_RAM_13 => X"0FFFFFFFFFFDB7FFF1FFFFF1FFFF7BDFF1999991F1DB7FF1F7777BDDFDDB7BDD",
            INIT_RAM_14 => X"FFFFF777F3D5B55BFFDB7F99F7173537F5BB1BB7FFFFFBBBF7F77777FFFFFFFF",
            INIT_RAM_15 => X"FFDB7FFFF7FFFFFFFFFF1FFFFB77FFFFFF77177FF7537357F7FFFFF7F7BDDDB7",
            INIT_RAM_16 => X"FBBB7FF1F3DD1DB7F3DFF1D1FFF1DB7FF3DF7FF1F1DB7FD3F3777737F3D95DD3",
            INIT_RAM_17 => X"F7F77FD3FB7FFF7BFFF1F1FFFF7BDB7FFB77F7FFFFF7F7FFF1FF3DD3F3DD3DD3",
            INIT_RAM_18 => X"F3DDDDD3FDDD1DD1F1DD1DD1F1DDDDD1F3DDDDD3F1DD1DD1FDD1DDB7F3D555D3",
            INIT_RAM_19 => X"F3DDDDD3FDDD59DDFDDD559DF1DDDDDDFDD595DDF3DFFFFFF3777773FDDD1DDD",
            INIT_RAM_1A => X"FD955DDDF7BDDDDDF3DDDDDDF7777771F3DF3DD3FDD51DD1F3D5DDD3FDDD1DD1",
            INIT_RAM_1B => X"0FFFFFFFFFFDB7FFF1FFFFF1FFFF7BDFF1999991F1DB7FF1F7777BDDFDDB7BDD",
            INIT_RAM_1C => X"3F3DD3FFFBBB1BB7F3D1D3FFF3DDD3FFF3DDD3FFF1DDD1DDF3D3F3FFFFFFFF7B",
            INIT_RAM_1D => X"F3DDD3FFFDDDD1FFFD5559FFF3777773FDD1DDDD3DFFF7FFF37773F7FDDDD1DD",
            INIT_RAM_1E => X"F955DDFFF7BDDDFFF3DDDDFFF7BBB1BBF1F3D3FFFDDD95FFFF3DD3FFDD1DD1FF",
            INIT_RAM_1F => X"FF5B5B5FFFFFFF53F177F77177777777F7339337F1B7F1FF3F3DDDFFFDB7BDFF",
            INIT_RAM_20 => X"FF882888FF996999FFAAAAAAFFBBEBBBFFCC3CCCFFDD7DDDFFEEBEEEFFFFFFFF",
            INIT_RAM_21 => X"FF000000FF114111FF228222FF33C333FF441444FF555555FF669666FF77D777",
            INIT_RAM_22 => X"BE882888BE996999BEAAAAAABEBBEBBBBECC3CCCBEDD7DDDBEEEBEEEBEFFFFFF",
            INIT_RAM_23 => X"BE000000BE114111BE228222BE33C333BE441444BE555555BE669666BE77D777",
            INIT_RAM_24 => X"7D8828887D9969997DAAAAAA7DBBEBBB7DCC3CCC7DDD7DDD7DEEBEEE7DFFFFFF",
            INIT_RAM_25 => X"7D0000007D1141117D2282227D33C3337D4414447D5555557D6696667D77D777",
            INIT_RAM_26 => X"3C8828883C9969993CAAAAAA3CBBEBBB3CCC3CCC3CDD7DDD3CEEBEEE3CFFFFFF",
            INIT_RAM_27 => X"3C0000003C1141113C2282223C33C3333C4414443C5555553C6696663C77D777",
            INIT_RAM_28 => X"EB882888EB996999EBAAAAAAEBBBEBBBEBCC3CCCEBDD7DDDEBEEBEEEEBFFFFFF",
            INIT_RAM_29 => X"EB000000EB114111EB228222EB33C333EB441444EB555555EB669666EB77D777",
            INIT_RAM_2A => X"AA882888AA996999AAAAAAAAAABBEBBBAACC3CCCAADD7DDDAAEEBEEEAAFFFFFF",
            INIT_RAM_2B => X"AA000000AA114111AA228222AA33C333AA441444AA555555AA669666AA77D777",
            INIT_RAM_2C => X"698828886999699969AAAAAA69BBEBBB69CC3CCC69DD7DDD69EEBEEE69FFFFFF",
            INIT_RAM_2D => X"6900000069114111692282226933C3336944144469555555696696666977D777",
            INIT_RAM_2E => X"288828882899699928AAAAAA28BBEBBB28CC3CCC28DD7DDD28EEBEEE28FFFFFF",
            INIT_RAM_2F => X"2800000028114111282282222833C3332844144428555555286696662877D777",
            INIT_RAM_30 => X"D7882888D7996999D7AAAAAAD7BBEBBBD7CC3CCCD7DD7DDDD7EEBEEED7FFFFFF",
            INIT_RAM_31 => X"D7000000D7114111D7228222D733C333D7441444D7555555D7669666D777D777",
            INIT_RAM_32 => X"968828889699699996AAAAAA96BBEBBB96CC3CCC96DD7DDD96EEBEEE96FFFFFF",
            INIT_RAM_33 => X"9600000096114111962282229633C3339644144496555555966696669677D777",
            INIT_RAM_34 => X"558828885599699955AAAAAA55BBEBBB55CC3CCC55DD7DDD55EEBEEE55FFFFFF",
            INIT_RAM_35 => X"5500000055114111552282225533C3335544144455555555556696665577D777",
            INIT_RAM_36 => X"148828881499699914AAAAAA14BBEBBB14CC3CCC14DD7DDD14EEBEEE14FFFFFF",
            INIT_RAM_37 => X"1400000014114111142282221433C3331444144414555555146696661477D777",
            INIT_RAM_38 => X"C3882888C3996999C3AAAAAAC3BBEBBBC3CC3CCCC3DD7DDDC3EEBEEEC3FFFFFF",
            INIT_RAM_39 => X"C3000000C3114111C3228222C333C333C3441444C3555555C3669666C377D777",
            INIT_RAM_3A => X"828828888299699982AAAAAA82BBEBBB82CC3CCC82DD7DDD82EEBEEE82FFFFFF",
            INIT_RAM_3B => X"8200000082114111822282228233C3338244144482555555826696668277D777",
            INIT_RAM_3C => X"418828884199699941AAAAAA41BBEBBB41CC3CCC41DD7DDD41EEBEEE41FFFFFF",
            INIT_RAM_3D => X"4100000041114111412282224133C3334144144441555555416696664177D777",
            INIT_RAM_3E => X"008828880099699900AAAAAA00BBEBBB00CC3CCC00DD7DDD00EEBEEE00FFFFFF",
            INIT_RAM_3F => X"0000000000114111002282220033C3330044144400555555006696660077D777"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 4,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0323000300001003030010030122222101200021012212210223221003013221",
            INIT_RAM_01 => X"0122222102232222022222320300000002100012012222220100000102223222",
            INIT_RAM_02 => X"0232222200122222012222220000000301221021021012210212222100001221",
            INIT_RAM_03 => X"7000000000021000033333330021000003000003030001230000012202210122",
            INIT_RAM_04 => X"0000000002120000033001200012103007000043000001110000000000000000",
            INIT_RAM_05 => X"0000012000000000000030000000000000003000002101200012221000000000",
            INIT_RAM_06 => X"0000012301221003012221030113111101221123030012210100000001222321",
            INIT_RAM_07 => X"0000012100012100000303000100000100000000000000000012322101221221",
            INIT_RAM_08 => X"8FFFFFEFFCC8C89888889AC8FFFFEDBF8DEFFED8BCEFFFFFCBDDBCFEC8CC8CFE",
            INIT_RAM_09 => X"9EEE8EEECCCCCCCCFF8BBBBBFFFFFFF8FFFFBDEFFEDBFFFFDFFFFFFFFFFF8FFF",
            INIT_RAM_0A => X"DADADADAADADADADFFED8DEF8FFFFFFFFFFF8FFFBBF8CEBBBBEC8FBB8FFECEF9",
            INIT_RAM_0B => X"FFFFFFFF8BBBBBB8FEE8F8EE8FFFFFF8FFEC8CEFBBBBBBBBF8BBBCFFF8FFFBCF",
            INIT_RAM_0C => X"1232210000001021030321000322232203000300012221000323210000000100",
            INIT_RAM_0D => X"0122210002222100022223000100000002101200011111010100000002222100",
            INIT_RAM_0E => X"0322220000122200023222000120010001210300000003002232230000122100",
            INIT_RAM_0F => X"0021212000000012001131100000000003000003030013001232220002101200",
            INIT_RAM_10 => X"FCDCFFFCFFFFEFFCFCFFEFFCFEDDDDDEFEDFFFDEFEDDEDDEFDDCDDEFFCFECDDE",
            INIT_RAM_11 => X"FEDDDDDEFDDCDDDDFDDDDDCDFCFFFFFFFDEFFFEDFEDDDDDDFEFFFFFEFDDDCDDD",
            INIT_RAM_12 => X"FDCDDDDDFFEDDDDDFEDDDDDDFFFFFFFCFEDDEFDEFDEFEDDEFDEDDDDEFFFFEDDE",
            INIT_RAM_13 => X"8FFFFFFFFFFDEFFFFCCCCCCCFFDEFFFFFCFFFFFCFCFFFEDCFFFFFEDDFDDEFEDD",
            INIT_RAM_14 => X"FFFFFFFFFDEDFFFFFCCFFEDFFFEDEFCFF8FFFFBCFFFFFEEEFFFFFFFFFFFFFFFF",
            INIT_RAM_15 => X"FFFFFEDFFFFFFFFFFFFFCFFFFFFFFFFFFFFFCFFFFFDEFEDFFFEDDDEFFFFFFFFF",
            INIT_RAM_16 => X"FFFFFEDCFEDDEFFCFEDDDEFCFEECEEEEFEDDEEDCFCFFEDDEFEFFFFFFFEDDDCDE",
            INIT_RAM_17 => X"FFFFFEDEFFFEDEFFFFFCFCFFFEFFFFFEFFFFFFFFFFFFFFFFFFEDCDDEFEDDEDDE",
            INIT_RAM_18 => X"FCDCFFFCFFFFEFFCFCFFEFFCFEDDDDDEFEDFFFDEFEDDEDDEFDDCDDEFFCFECDDE",
            INIT_RAM_19 => X"FEDDDDDEFDDCDDDDFDDDDDCDFCFFFFFFFDEFFFEDFEDDDDDDFEFFFFFEFDDDCDDD",
            INIT_RAM_1A => X"FDCDDDDDFFEDDDDDFEDDDDDDFFFFFFFCFEDDEFDEFDEFEDDEFDEDDDDEFFFFEDDE",
            INIT_RAM_1B => X"8FFFFFFFFFFDEFFFFCCCCCCCFFDEFFFFFCFFFFFCFCFFFEDCFFFFFEDDFDDEFEDD",
            INIT_RAM_1C => X"EDCDDEFFFFFFEFDEFCFCDEFFFCDDDCDDFCFFFCFFFEDDDEFFFCDCDEFFFFFFFEFF",
            INIT_RAM_1D => X"FEDDDEFFFDDDDEFFFDDDDCFFFEFFFFFFFDEFEDFFFEEEEEFEFEFFFFFFFDDDDEFF",
            INIT_RAM_1E => X"FCDDDDFFFFEDDDFFFDCDDDFFFEDFFEFFFEDEFCFFFFFFFCFFDDCDDCFFFFEDDEFF",
            INIT_RAM_1F => X"FFDEDEDFFFFFFFEDFFEECEEFFFFFFFFFFCFFFFFCFCFFECFFEDCDDDFFFDEFEDFF",
            INIT_RAM_20 => X"FFFF28FFFFFF69FFFFFFAAFFFFFFEBFFFFFF3CFFFFFF7DFFFFFFBEFFFFFFFFFF",
            INIT_RAM_21 => X"FFFF00FFFFFF41FFFFFF82FFFFFFC3FFFFFF14FFFFFF55FFFFFF96FFFFFFD7FF",
            INIT_RAM_22 => X"BEEE28EEBEEE69EEBEEEAAEEBEEEEBEEBEEE3CEEBEEE7DEEBEEEBEEEBEEEFFEE",
            INIT_RAM_23 => X"BEEE00EEBEEE41EEBEEE82EEBEEEC3EEBEEE14EEBEEE55EEBEEE96EEBEEED7EE",
            INIT_RAM_24 => X"7DDD28DD7DDD69DD7DDDAADD7DDDEBDD7DDD3CDD7DDD7DDD7DDDBEDD7DDDFFDD",
            INIT_RAM_25 => X"7DDD00DD7DDD41DD7DDD82DD7DDDC3DD7DDD14DD7DDD55DD7DDD96DD7DDDD7DD",
            INIT_RAM_26 => X"3CCC28CC3CCC69CC3CCCAACC3CCCEBCC3CCC3CCC3CCC7DCC3CCCBECC3CCCFFCC",
            INIT_RAM_27 => X"3CCC00CC3CCC41CC3CCC82CC3CCCC3CC3CCC14CC3CCC55CC3CCC96CC3CCCD7CC",
            INIT_RAM_28 => X"EBBB28BBEBBB69BBEBBBAABBEBBBEBBBEBBB3CBBEBBB7DBBEBBBBEBBEBBBFFBB",
            INIT_RAM_29 => X"EBBB00BBEBBB41BBEBBB82BBEBBBC3BBEBBB14BBEBBB55BBEBBB96BBEBBBD7BB",
            INIT_RAM_2A => X"AAAA28AAAAAA69AAAAAAAAAAAAAAEBAAAAAA3CAAAAAA7DAAAAAABEAAAAAAFFAA",
            INIT_RAM_2B => X"AAAA00AAAAAA41AAAAAA82AAAAAAC3AAAAAA14AAAAAA55AAAAAA96AAAAAAD7AA",
            INIT_RAM_2C => X"69992899699969996999AA996999EB9969993C9969997D996999BE996999FF99",
            INIT_RAM_2D => X"6999009969994199699982996999C3996999149969995599699996996999D799",
            INIT_RAM_2E => X"28882888288869882888AA882888EB8828883C8828887D882888BE882888FF88",
            INIT_RAM_2F => X"2888008828884188288882882888C3882888148828885588288896882888D788",
            INIT_RAM_30 => X"D7FF28FFD7FF69FFD7FFAAFFD7FFEBFFD7FF3CFFD7FF7DFFD7FFBEFFD7FFFFFF",
            INIT_RAM_31 => X"D7FF00FFD7FF41FFD7FF82FFD7FFC3FFD7FF14FFD7FF55FFD7FF96FFD7FFD7FF",
            INIT_RAM_32 => X"96EE28EE96EE69EE96EEAAEE96EEEBEE96EE3CEE96EE7DEE96EEBEEE96EEFFEE",
            INIT_RAM_33 => X"96EE00EE96EE41EE96EE82EE96EEC3EE96EE14EE96EE55EE96EE96EE96EED7EE",
            INIT_RAM_34 => X"55DD28DD55DD69DD55DDAADD55DDEBDD55DD3CDD55DD7DDD55DDBEDD55DDFFDD",
            INIT_RAM_35 => X"55DD00DD55DD41DD55DD82DD55DDC3DD55DD14DD55DD55DD55DD96DD55DDD7DD",
            INIT_RAM_36 => X"14CC28CC14CC69CC14CCAACC14CCEBCC14CC3CCC14CC7DCC14CCBECC14CCFFCC",
            INIT_RAM_37 => X"14CC00CC14CC41CC14CC82CC14CCC3CC14CC14CC14CC55CC14CC96CC14CCD7CC",
            INIT_RAM_38 => X"C3BB28BBC3BB69BBC3BBAABBC3BBEBBBC3BB3CBBC3BB7DBBC3BBBEBBC3BBFFBB",
            INIT_RAM_39 => X"C3BB00BBC3BB41BBC3BB82BBC3BBC3BBC3BB14BBC3BB55BBC3BB96BBC3BBD7BB",
            INIT_RAM_3A => X"82AA28AA82AA69AA82AAAAAA82AAEBAA82AA3CAA82AA7DAA82AABEAA82AAFFAA",
            INIT_RAM_3B => X"82AA00AA82AA41AA82AA82AA82AAC3AA82AA14AA82AA55AA82AA96AA82AAD7AA",
            INIT_RAM_3C => X"41992899419969994199AA994199EB9941993C9941997D994199BE994199FF99",
            INIT_RAM_3D => X"4199009941994199419982994199C3994199149941995599419996994199D799",
            INIT_RAM_3E => X"00882888008869880088AA880088EB8800883C8800887D880088BE880088FF88",
            INIT_RAM_3F => X"0088008800884188008882880088C3880088148800885588008896880088D788"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

end Behavioral; --Gowin_pROM_video
