--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.10.03 (64-bit)
--Part Number: GW5AT-LV60PG484AC1/I0
--Device: GW5AT-60
--Device Version: B
--Created Time: Wed May 28 16:04:34 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_key is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(10 downto 0)
    );
end Gowin_pROM_key;

architecture Behavioral of Gowin_pROM_key is

    signal prom_inst_0_dout_w: std_logic_vector(23 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dout(7 downto 0) <= prom_inst_0_DO_o(7 downto 0) ;
    prom_inst_0_dout_w(23 downto 0) <= prom_inst_0_DO_o(31 downto 8) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 8,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"3726372635253525365E1E1E342434243323332332400000312131211B1B1B1B",
            INIT_RAM_01 => X"59591919525212124545050557571717515111110909090939283928382A382A",
            INIT_RAM_02 => X"484808085353131344440404414101014F4F0F0F494909095555151554541414",
            INIT_RAM_03 => X"585818185A5A1A1A4C4C0C0C3B3A3B3A4B4B0B0B4A4A0A0A4747070746460606",
            INIT_RAM_04 => X"2F3F2F3F2E3E2E3E2C3C2C3C4D4D0D0D4E4E0E0E424202025656161643430303",
            INIT_RAM_05 => X"3D2B3D2B607E607E33333333323232323131313130303030080808082F2F2F2F",
            INIT_RAM_06 => X"373737373636363635353535343434341B1B1B1B292929292D5F1F1F30293029",
            INIT_RAM_07 => X"3939393938383838151515152A2A2A2A5D7D1D1D5B7B1B1B505010105C7C1C1C",
            INIT_RAM_08 => X"202020203F3F3F3F27222722202020200B0B0B0B0D0D0D0D2B2B2B2B2E2E2E2E",
            INIT_RAM_09 => X"15151515080808080A0A0A0A7F7F7F7F2C2C2C2C0D0D0D0D2D2D2D2D28282828",
            INIT_RAM_0A => X"204120204D20202020202020202020202020204E20204820204F20204A202020",
            INIT_RAM_0B => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A02020204420204320",
            INIT_RAM_0C => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_0D => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_0E => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_0F => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_10 => X"3726372635253525365E1E1E342434243323332332400000312131211B1B1B1B",
            INIT_RAM_11 => X"79591919725212126545050577571717715111110909090939283928382A382A",
            INIT_RAM_12 => X"684808087353131364440404614101016F4F0F0F694909097555151574541414",
            INIT_RAM_13 => X"785818187A5A1A1A6C4C0C0C3B3A3B3A6B4B0B0B6A4A0A0A6747070766460606",
            INIT_RAM_14 => X"2F3F2F3F2E3E2E3E2C3C2C3C6D4D0D0D6E4E0E0E624202027656161663430303",
            INIT_RAM_15 => X"3D2B3D2B607E607E33333333323232323131313130303030080808082F2F2F2F",
            INIT_RAM_16 => X"373737373636363635353535343434341B1B1B1B292929292D5F1F1F30293029",
            INIT_RAM_17 => X"3939393938383838151515152A2A2A2A5D7D1D1D5B7B1B1B705010105C7C1C1C",
            INIT_RAM_18 => X"202020203F3F3F3F27222722202020200B0B0B0B0D0D0D0D2B2B2B2B2E2E2E2E",
            INIT_RAM_19 => X"15151515080808080A0A0A0A7F7F7F7F2C2C2C2C0D0D0D0D2D2D2D2D28282828",
            INIT_RAM_1A => X"204120204D20202020202020202020202020204E20204820204F20204A202020",
            INIT_RAM_1B => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A02020204420204320",
            INIT_RAM_1C => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_1D => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_1E => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_1F => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_20 => X"3726372635253525365E1E1E342434243323332332400000312131211B1B1B1B",
            INIT_RAM_21 => X"59591919525212124545050557571717515111110909090939283928382A382A",
            INIT_RAM_22 => X"484808085353131344440404414101014F4F0F0F494909095555151554541414",
            INIT_RAM_23 => X"585818185A5A1A1A4C4C0C0C3B3A3B3A4B4B0B0B4A4A0A0A4747070746460606",
            INIT_RAM_24 => X"2F3F2F3F2E3E2E3E2C3C2C3C4D4D0D0D4E4E0E0E424202025656161643430303",
            INIT_RAM_25 => X"3D2B3D2B607E607E33333333323232323131313130303030080808082F2F2F2F",
            INIT_RAM_26 => X"373737373636363635353535343434341B1B1B1B292929292D5F1F1F30293029",
            INIT_RAM_27 => X"3939393938383838151515152A2A2A2A5D7D1D1D5B7B1B1B505010105C7C1C1C",
            INIT_RAM_28 => X"202020203F3F3F3F27222722202020200B0B0B0B0D0D0D0D2B2B2B2B2E2E2E2E",
            INIT_RAM_29 => X"15151515080808080A0A0A0A7F7F7F7F2C2C2C2C0D0D0D0D2D2D2D2D28282828",
            INIT_RAM_2A => X"204120204D20202020202020202020202020204E20204820204F20204A202020",
            INIT_RAM_2B => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A02020204420204320",
            INIT_RAM_2C => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_2D => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_2E => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_2F => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_30 => X"3726372635253525365E1E1E342434243323332332400000312131211B1B1B1B",
            INIT_RAM_31 => X"79591919725212126545050577571717715111110909090939283928382A382A",
            INIT_RAM_32 => X"684808087353131364440404614101016F4F0F0F694909097555151574541414",
            INIT_RAM_33 => X"785818187A5A1A1A6C4C0C0C3B3A3B3A6B4B0B0B6A4A0A0A6747070766460606",
            INIT_RAM_34 => X"2F3F2F3F2E3E2E3E2C3C2C3C6D4D0D0D6E4E0E0E624202027656161663430303",
            INIT_RAM_35 => X"3D2B3D2B607E607E33333333323232323131313130303030080808082F2F2F2F",
            INIT_RAM_36 => X"373737373636363635353535343434341B1B1B1B292929292D5F1F1F30293029",
            INIT_RAM_37 => X"3939393938383838151515152A2A2A2A5D7D1D1D5B7B1B1B705010105C7C1C1C",
            INIT_RAM_38 => X"202020203F3F3F3F27222722202020200B0B0B0B0D0D0D0D2B2B2B2B2E2E2E2E",
            INIT_RAM_39 => X"15151515080808080A0A0A0A7F7F7F7F2C2C2C2C0D0D0D0D2D2D2D2D28282828",
            INIT_RAM_3A => X"204120204D20202020202020202020202020204E20204820204F20204A202020",
            INIT_RAM_3B => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A02020204420204320",
            INIT_RAM_3C => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_3D => X"A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_3E => X"303531302D313433A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0",
            INIT_RAM_3F => X"32383931A052455455504D4F43A0454C505041A0544847495259504F43A0A041"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

end Behavioral; --Gowin_pROM_key
