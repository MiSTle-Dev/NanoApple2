
module Gowin_pROM_uc (dout, clk, oce, ce, reset, ad);

output [39:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [26:0] promx9_inst_0_dout_w;
wire [8:0] promx9_inst_0_dout;
wire [26:0] promx9_inst_1_dout_w;
wire [8:0] promx9_inst_1_dout;
wire [26:0] promx9_inst_2_dout_w;
wire [17:9] promx9_inst_2_dout;
wire [26:0] promx9_inst_3_dout_w;
wire [17:9] promx9_inst_3_dout;
wire [26:0] promx9_inst_4_dout_w;
wire [26:18] promx9_inst_4_dout;
wire [26:0] promx9_inst_5_dout_w;
wire [26:18] promx9_inst_5_dout;
wire [26:0] promx9_inst_6_dout_w;
wire [35:27] promx9_inst_6_dout;
wire [26:0] promx9_inst_7_dout_w;
wire [35:27] promx9_inst_7_dout;
wire [27:0] prom_inst_8_dout_w;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[11])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[11])
);
defparam lut_inst_1.INIT = 4'h8;
pROMX9 promx9_inst_0 (
    .DO({promx9_inst_0_dout_w[26:0],promx9_inst_0_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_0.READ_MODE = 1'b0;
defparam promx9_inst_0.BIT_WIDTH = 9;
defparam promx9_inst_0.RESET_MODE = "SYNC";
defparam promx9_inst_0.INIT_RAM_00 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_01 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_02 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_03 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_04 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_05 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_06 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_07 = 288'h000000000000008200080000600000000000000000000000010200080000800000000000;
defparam promx9_inst_0.INIT_RAM_08 = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_09 = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_0A = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_0B = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_0C = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_0D = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_0E = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_0F = 288'h000000000000000600000000000000000000000000000000000800000000000000000000;
defparam promx9_inst_0.INIT_RAM_10 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_11 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_12 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_13 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_14 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_15 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_16 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_17 = 288'h000000000000000000000440010000000020000000000000000000000440010000000020;
defparam promx9_inst_0.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000200000000000000000000;
defparam promx9_inst_0.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000E00000000000000000000;
defparam promx9_inst_0.INIT_RAM_1B = 288'h000000000000000E00000000000000000000000000000000020E00000000000000000000;
defparam promx9_inst_0.INIT_RAM_1C = 288'h000000000000020C00000000000000000000000000000000000C00000000000000000000;
defparam promx9_inst_0.INIT_RAM_1D = 288'h000000000000000000000000000000240000000000000000001200000000000000000000;
defparam promx9_inst_0.INIT_RAM_1E = 288'h000000000000000000000001200000000000000000000000000200000000000000000000;
defparam promx9_inst_0.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000008000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000038000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_23 = 288'h000000000038000000000000000000000000000000000838000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_24 = 288'h000000000830000000000000000000000000000000000030000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_25 = 288'h000000000000000000000000009000240000000000000048000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_26 = 288'h000000000048000000000000000000000000000000000008000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000008000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000038000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_2B = 288'h000000000038000000000000000000000000000000000838000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_2C = 288'h000000000830000000000000000000000000000000000030000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000048000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_2E = 288'h000000000048000000000000000000000000000000000008000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000001000000000000000000;
defparam promx9_inst_0.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000007000000000000000000;
defparam promx9_inst_0.INIT_RAM_33 = 288'h000000000000000007000000000000000000000000000000000107000000000000000000;
defparam promx9_inst_0.INIT_RAM_34 = 288'h000000000000000106000000000000000000000000000000000006000000000000000000;
defparam promx9_inst_0.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000009000000000000000000;
defparam promx9_inst_0.INIT_RAM_36 = 288'h000000000000000000000000009000000000000000000000000001000000000000000000;
defparam promx9_inst_0.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000040000000000000000000000;
defparam promx9_inst_0.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_3A = 288'h0000000000000000000000000000000000000000000000001C0000000000000000000000;
defparam promx9_inst_0.INIT_RAM_3B = 288'h0000000000001C00000000000000000000000000000000041C0000000000000000000000;
defparam promx9_inst_0.INIT_RAM_3C = 288'h000000000004180000000000000000000000000000000000180000000000000000000000;
defparam promx9_inst_0.INIT_RAM_3D = 288'h000000000000000200000040000008000200000000000000240000000000000000000000;
defparam promx9_inst_0.INIT_RAM_3E = 288'h000000000000000000000240000000000000000000000000040000000000000000000000;
defparam promx9_inst_0.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

pROMX9 promx9_inst_1 (
    .DO({promx9_inst_1_dout_w[26:0],promx9_inst_1_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_1.READ_MODE = 1'b0;
defparam promx9_inst_1.BIT_WIDTH = 9;
defparam promx9_inst_1.RESET_MODE = "SYNC";
defparam promx9_inst_1.INIT_RAM_00 = 288'h000000000000000000000000200008000000000000000000000000000000001000000000;
defparam promx9_inst_1.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000008000000;
defparam promx9_inst_1.INIT_RAM_02 = 288'h000000000000000000000000200000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_0A = 288'h000000000000000000008000000000000000000000000000000000008000000000000000;
defparam promx9_inst_1.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000008000000000000000;
defparam promx9_inst_1.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_10 = 288'h000000000000000000000240000000000000000000000000000000000240000000000000;
defparam promx9_inst_1.INIT_RAM_11 = 288'h000000000000000000000240000000000000000000000000000000004240000000000000;
defparam promx9_inst_1.INIT_RAM_12 = 288'h000000000000000000000080000000000000000000000000000000000080000000000000;
defparam promx9_inst_1.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_14 = 288'h000000000000000000004040000000000000000000000000000000000140000000000000;
defparam promx9_inst_1.INIT_RAM_15 = 288'h000000000000000000000040000000000000000000000000000000000200000000000000;
defparam promx9_inst_1.INIT_RAM_16 = 288'h000000000000000000000040010000040000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_18 = 288'h000000000000000000000240000000000000000000000000000000000240000000000000;
defparam promx9_inst_1.INIT_RAM_19 = 288'h000000000000000000000240000000000000000000000000000000004240000000000000;
defparam promx9_inst_1.INIT_RAM_1A = 288'h000000000000000000000080000000000000000000000000000000000080000000000000;
defparam promx9_inst_1.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_1C = 288'h000000000000000000004040000000000000000000000000000000000140000000000000;
defparam promx9_inst_1.INIT_RAM_1D = 288'h000000000000000000000040000000000000000000000000000000000200000000000000;
defparam promx9_inst_1.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_20 = 288'h000000000000000000000001200000000000000000000000000000000001200000000000;
defparam promx9_inst_1.INIT_RAM_21 = 288'h000000000000000000000001200000000000000000000000000000000021200000000000;
defparam promx9_inst_1.INIT_RAM_22 = 288'h000000000000000000000000400000000000000000000000000000000000400000000000;
defparam promx9_inst_1.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_24 = 288'h000000000000000000000020200000000000000000000000000000000000A00000000000;
defparam promx9_inst_1.INIT_RAM_25 = 288'h000000000000000000000000200000000000000000000000000000000001000000000000;
defparam promx9_inst_1.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_28 = 288'h000000000000001200000000000000000000000000000000001200000000000000000000;
defparam promx9_inst_1.INIT_RAM_29 = 288'h000000000000001200000000000000000000000000000000021200000000000000000000;
defparam promx9_inst_1.INIT_RAM_2A = 288'h000000000000000400000000000000000000000000000000000400000000000000000000;
defparam promx9_inst_1.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_2C = 288'h000000000000020200000000000000000000000000000000000A00000000000000000000;
defparam promx9_inst_1.INIT_RAM_2D = 288'h000000000000000200000000000000000000000000000000001000000000000000000000;
defparam promx9_inst_1.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_30 = 288'h000000000000000000000001200000000000000000000000000000000001200000000000;
defparam promx9_inst_1.INIT_RAM_31 = 288'h000000000000000000000001200000000000000000000000000000000021200000000000;
defparam promx9_inst_1.INIT_RAM_32 = 288'h000000000000000000000000400000000000000000000000000000000000400000000000;
defparam promx9_inst_1.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_34 = 288'h000000000000000000000020200000000000000000000000000000000000A00000000000;
defparam promx9_inst_1.INIT_RAM_35 = 288'h000000000000000000000000200000000000000000000000000000000001000000000000;
defparam promx9_inst_1.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_38 = 288'h000000000000000000048000000000000000000000000000000000048000000000000000;
defparam promx9_inst_1.INIT_RAM_39 = 288'h000000000000000000048000000000000000000000000000000000848000000000000000;
defparam promx9_inst_1.INIT_RAM_3A = 288'h000000000000000000010000000000000000000000000000000000010000000000000000;
defparam promx9_inst_1.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_3C = 288'h000000000000000000808000000000000000000000000000000000028000000000000000;
defparam promx9_inst_1.INIT_RAM_3D = 288'h000000000000000000008000000000000000000000000000000000040000000000000000;
defparam promx9_inst_1.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_1.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

pROMX9 promx9_inst_2 (
    .DO({promx9_inst_2_dout_w[26:0],promx9_inst_2_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_2.READ_MODE = 1'b0;
defparam promx9_inst_2.BIT_WIDTH = 9;
defparam promx9_inst_2.RESET_MODE = "SYNC";
defparam promx9_inst_2.INIT_RAM_00 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_01 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_02 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_03 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_04 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_05 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_06 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_07 = 288'h000000000800000000000000400000000000000000000800000000000000400000000000;
defparam promx9_inst_2.INIT_RAM_08 = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_09 = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_0A = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_0B = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_0C = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_0D = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_0E = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_0F = 288'h000000100001000000000000000000000000000000100001000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_10 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_11 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_12 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_13 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_14 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_15 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_16 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_17 = 288'h000000000000000100000000000000000000000000000000000100000000000000000000;
defparam promx9_inst_2.INIT_RAM_18 = 288'h00000000000000000000000000000000002C000000100001002400000000000000000000;
defparam promx9_inst_2.INIT_RAM_19 = 288'h00000010000100280000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_1A = 288'h00000000000000000000000000000000002C000000100001002400000000000000000000;
defparam promx9_inst_2.INIT_RAM_1B = 288'h000000100001002600000000000000000000000000100001002400000000000000000000;
defparam promx9_inst_2.INIT_RAM_1C = 288'h000000100001002400000000000000000000000000100001002400000000000000000000;
defparam promx9_inst_2.INIT_RAM_1D = 288'h000000000000000000000000000001000000000000100001002000000000000000000000;
defparam promx9_inst_2.INIT_RAM_1E = 288'h000000000000000100001002000000000000000000100001002000000000000000000000;
defparam promx9_inst_2.INIT_RAM_1F = 288'h000000100001001C0000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_20 = 288'h00000000000000000000000000000000002C000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_21 = 288'h0000000000A400000000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_22 = 288'h00000000000000000000000000000000002C000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_23 = 288'h00000000009C000000000000000000000000000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_24 = 288'h000000000094000000000000000000000000000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_25 = 288'h000000000000000000000000080402010080000000000084000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_26 = 288'h000000000084000000000000000000000000000000000084000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_27 = 288'h00000000007400000000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_28 = 288'h00000000000000000000000000000000002C000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_29 = 288'h0000000000A400000000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_2A = 288'h00000000000000000000000000000000002C000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_2B = 288'h00000000009C000000000000000000000000000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_2C = 288'h000000000094000000000000000000000000000000000094000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_2D = 288'h00000000000000000000000000000000002C000000000084000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_2E = 288'h000000000084000000000000000000000000000000000084000000000000000000000000;
defparam promx9_inst_2.INIT_RAM_2F = 288'h00000000007400000000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_30 = 288'h00000000000000000000000000000000002C000000000800008012000000000000000000;
defparam promx9_inst_2.INIT_RAM_31 = 288'h00000000080000801400000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_32 = 288'h00000000000000000000000000000000002C000000000800008012000000000000000000;
defparam promx9_inst_2.INIT_RAM_33 = 288'h000000000800008013000000000000000000000000000800008012000000000000000000;
defparam promx9_inst_2.INIT_RAM_34 = 288'h000000000800008012000000000000000000000000000800008012000000000000000000;
defparam promx9_inst_2.INIT_RAM_35 = 288'h00000000000000000000000000000000002C000000000800008010000000000000000000;
defparam promx9_inst_2.INIT_RAM_36 = 288'h000000000000000000800008010000000000000000000800008010000000000000000000;
defparam promx9_inst_2.INIT_RAM_37 = 288'h00000000080000800E00000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_38 = 288'h00000000000000000000000000000000002C000020000200480000000000000000000000;
defparam promx9_inst_2.INIT_RAM_39 = 288'h00002000020050000000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_2.INIT_RAM_3A = 288'h00000000000000000000000000000000002C000020000200480000000000000000000000;
defparam promx9_inst_2.INIT_RAM_3B = 288'h0000200002004C0000000000000000000000000020000200480000000000000000000000;
defparam promx9_inst_2.INIT_RAM_3C = 288'h000020000200480000000000000000000000000020000200480000000000000000000000;
defparam promx9_inst_2.INIT_RAM_3D = 288'h000000000402030080406010080C02000000000020000200400000000000000000000000;
defparam promx9_inst_2.INIT_RAM_3E = 288'h000000000000020000200400000000000000000020000200400000000000000000000000;
defparam promx9_inst_2.INIT_RAM_3F = 288'h00002000020038000000000000000000000000000000000000000000000000000000002C;

pROMX9 promx9_inst_3 (
    .DO({promx9_inst_3_dout_w[26:0],promx9_inst_3_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_3.READ_MODE = 1'b0;
defparam promx9_inst_3.BIT_WIDTH = 9;
defparam promx9_inst_3.RESET_MODE = "SYNC";
defparam promx9_inst_3.INIT_RAM_00 = 288'h000000000000020000006030080000000000000000000000020080006010180000000000;
defparam promx9_inst_3.INIT_RAM_01 = 288'h00001008040201008040000000000000008C00000000000000010C000028040A01000000;
defparam promx9_inst_3.INIT_RAM_02 = 288'h000000000000000000000000000000020000000000000000000000000000000004000100;
defparam promx9_inst_3.INIT_RAM_03 = 288'h00000000000000000000000000000000010000000000000000000000000000000000002C;
defparam promx9_inst_3.INIT_RAM_04 = 288'h00000000000000000000000000000000002C00000000000000000000000000000000002C;
defparam promx9_inst_3.INIT_RAM_05 = 288'h00000000000000000000000000000000002C00000000000000000000000000000000002C;
defparam promx9_inst_3.INIT_RAM_06 = 288'h00000000000000000000000000000000002C00000000000000000000000000000000002C;
defparam promx9_inst_3.INIT_RAM_07 = 288'h00000000000000000010000000000000000A00000000000000000010000000000000000A;
defparam promx9_inst_3.INIT_RAM_08 = 288'h000000000000000000000000140200000100000000000000000000000000000000000100;
defparam promx9_inst_3.INIT_RAM_09 = 288'h000000000000000000000000000A01000000000000000000028040000000000004000100;
defparam promx9_inst_3.INIT_RAM_0A = 288'h000000000000028040000000000800020000000000000000028040000000000000020000;
defparam promx9_inst_3.INIT_RAM_0B = 288'h000000000000000000004000000000000000000000000000000000000000000800020000;
defparam promx9_inst_3.INIT_RAM_0C = 288'h000000000000000000034000000000000000000000000000000000024000000000000000;
defparam promx9_inst_3.INIT_RAM_0D = 288'h000000000000000000064000000000000000000000000000000000054000000000000000;
defparam promx9_inst_3.INIT_RAM_0E = 288'h000000000000000000004000000000000000000000000000000000004000000000000000;
defparam promx9_inst_3.INIT_RAM_0F = 288'h000000000000000000004000000000000000000000000002010080402010080000000080;
defparam promx9_inst_3.INIT_RAM_10 = 288'h0000000000000000000004A00000000000000000000000000000000004A0000000000000;
defparam promx9_inst_3.INIT_RAM_11 = 288'h0000000000000000000004A00000000000000000000000000000000004A0000000000000;
defparam promx9_inst_3.INIT_RAM_12 = 288'h000000000000000000000420000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_13 = 288'h00000000000000000000000000000000002C000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_14 = 288'h000000000000000000000220000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_15 = 288'h000000000000000000000220000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_16 = 288'h00000000000002000000000000000000000000000000000000000000000000000000002C;
defparam promx9_inst_3.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_18 = 288'h0000000000000000000004A00000000000000000000000000000000004A0000000000000;
defparam promx9_inst_3.INIT_RAM_19 = 288'h0000000000000000000004A00000000000000000000000000000000004A0000000000000;
defparam promx9_inst_3.INIT_RAM_1A = 288'h000000000000000000000420000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_1B = 288'h000000000004008010000000000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_1C = 288'h000000000000000000000220000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_1D = 288'h000000000000000000000220000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_1E = 288'h000000000000020000000000000000000000000000000000000000000000000004000000;
defparam promx9_inst_3.INIT_RAM_1F = 288'h000000000004008010000000000000000000000000000000000000000420000000000000;
defparam promx9_inst_3.INIT_RAM_20 = 288'h000000000000000000000002500000000000000000000000000000000002500000000000;
defparam promx9_inst_3.INIT_RAM_21 = 288'h000000000000000000000002500000000000000000000000000000000002500000000000;
defparam promx9_inst_3.INIT_RAM_22 = 288'h000000000000000000000002100000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_23 = 288'h000000000801002000000000000000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_24 = 288'h000000000000000000000001100000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_25 = 288'h000000000000000000000001100000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_26 = 288'h000000000004000000000000000000000000000000000000000000000000000800000000;
defparam promx9_inst_3.INIT_RAM_27 = 288'h000000000801002000000000000000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_28 = 288'h000000000000002500000000000000000000000000000000002500000000000000000000;
defparam promx9_inst_3.INIT_RAM_29 = 288'h000000000000002500000000000000000000000000000000002500000000000000000000;
defparam promx9_inst_3.INIT_RAM_2A = 288'h000000000000002100000000000000000000000000000000002100000000000000000000;
defparam promx9_inst_3.INIT_RAM_2B = 288'h000020040080000000000000000000000000000000000000002100000000000000000000;
defparam promx9_inst_3.INIT_RAM_2C = 288'h000000000000001100000000000000000000000000000000002100000000000000000000;
defparam promx9_inst_3.INIT_RAM_2D = 288'h000000000000001100000000000000000000000000000000002100000000000000000000;
defparam promx9_inst_3.INIT_RAM_2E = 288'h000000100000000000000000000000000000000000000000000000000020000000000000;
defparam promx9_inst_3.INIT_RAM_2F = 288'h000020040080000000000000000000000000000000000000002100000000000000000000;
defparam promx9_inst_3.INIT_RAM_30 = 288'h000000000000000000000002500000000000000000000000000000000002500000000000;
defparam promx9_inst_3.INIT_RAM_31 = 288'h000000000000000000000002500000000000000000000000000000000002500000000000;
defparam promx9_inst_3.INIT_RAM_32 = 288'h000000000000000000000002100000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_33 = 288'h000000000801002000000000000000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_34 = 288'h000000000000000000000001100000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_35 = 288'h000000000000000000000001100000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_36 = 288'h000000000004000000000000000000000000000000000000000000000000000800000000;
defparam promx9_inst_3.INIT_RAM_37 = 288'h000000000801002000000000000000000000000000000000000000000002100000000000;
defparam promx9_inst_3.INIT_RAM_38 = 288'h000000000000000000094000000000000000000000000000000000094000000000000000;
defparam promx9_inst_3.INIT_RAM_39 = 288'h000000000000000000094000000000000000000000000000000000094000000000000000;
defparam promx9_inst_3.INIT_RAM_3A = 288'h000000000000000000084000000000000000000000000000000000084000000000000000;
defparam promx9_inst_3.INIT_RAM_3B = 288'h000020040080000000000000000000000000000000000000000000084000000000000000;
defparam promx9_inst_3.INIT_RAM_3C = 288'h000000000000000000044000000000000000000000000000000000084000000000000000;
defparam promx9_inst_3.INIT_RAM_3D = 288'h000000000000000000044000000000000000000000000000000000084000000000000000;
defparam promx9_inst_3.INIT_RAM_3E = 288'h000000100000000000000000000000000000000000000000000000000020000000000000;
defparam promx9_inst_3.INIT_RAM_3F = 288'h000020040080000000000000000000000000000000000000000000084000000000000000;

pROMX9 promx9_inst_4 (
    .DO({promx9_inst_4_dout_w[26:0],promx9_inst_4_dout[26:18]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_4.READ_MODE = 1'b0;
defparam promx9_inst_4.BIT_WIDTH = 9;
defparam promx9_inst_4.RESET_MODE = "SYNC";
defparam promx9_inst_4.INIT_RAM_00 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_01 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_02 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_03 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_04 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_05 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_06 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_07 = 288'h0000200000000140000002C00000080000000000200000000140000002C0000008000000;
defparam promx9_inst_4.INIT_RAM_08 = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_09 = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_0A = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_0B = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_0C = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_0D = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_0E = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_0F = 288'h004000000000010000008000000000000000004000000000010000008000000000000000;
defparam promx9_inst_4.INIT_RAM_10 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_11 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_12 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_13 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_14 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_15 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_16 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_17 = 288'h00000000000400000000280000000000000B00000000000400000000280000000000000B;
defparam promx9_inst_4.INIT_RAM_18 = 288'h000000000000000000000000000000000000004000000000010000000000000000000001;
defparam promx9_inst_4.INIT_RAM_19 = 288'h004000000000010000000000000000000001000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_1A = 288'h000000000000000000000000000000000000004000000000010000000000000000000001;
defparam promx9_inst_4.INIT_RAM_1B = 288'h004000000000010000000000000000000001004000000000010000000000000000000001;
defparam promx9_inst_4.INIT_RAM_1C = 288'h004000000000010000000000000000000001004000000000010000000000000000000001;
defparam promx9_inst_4.INIT_RAM_1D = 288'h0000000000000000000000000000033CC000004000000000010000000000000000000001;
defparam promx9_inst_4.INIT_RAM_1E = 288'h000000000004000000000010000000000001004000000000010000000000000000000001;
defparam promx9_inst_4.INIT_RAM_1F = 288'h004000000000010000000000000000000001000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000900000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_21 = 288'h000000000900000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000900000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_23 = 288'h000000000900000000000000000000000000000000000900000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_24 = 288'h000000000900000000000000000000000000000000000900000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_25 = 288'h0000000000000000000000000CF003000000000000000900000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_26 = 288'h000000000800000000000000000000000000000000000900000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_27 = 288'h000000000900000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000F00000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_29 = 288'h000000000F00000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000F00000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_2B = 288'h000000000F00000000000000000000000000000000000F00000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_2C = 288'h000000000F00000000000000000000000000000000000F00000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000F00000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_2E = 288'h000000000800000000000000000000000000000000000F00000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_2F = 288'h000000000F00000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_30 = 288'h000000000000000000000000000000000000000020000000000080000000000000000009;
defparam promx9_inst_4.INIT_RAM_31 = 288'h000020000000000080000000000000000009000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_32 = 288'h000000000000000000000000000000000000000020000000000080000000000000000009;
defparam promx9_inst_4.INIT_RAM_33 = 288'h000020000000000080000000000000000009000020000000000080000000000000000009;
defparam promx9_inst_4.INIT_RAM_34 = 288'h000020000000000080000000000000000009000020000000000080000000000000000009;
defparam promx9_inst_4.INIT_RAM_35 = 288'h000000000000000000000000000000000000000020000000000080000000000000000009;
defparam promx9_inst_4.INIT_RAM_36 = 288'h000000000000020000000000080000000009000020000000000080000000000000000009;
defparam promx9_inst_4.INIT_RAM_37 = 288'h000020000000000080000000000000000009000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_38 = 288'h000000000000000000000000000000000000800000000002000000000000000000000006;
defparam promx9_inst_4.INIT_RAM_39 = 288'h800000000002000000000000000000000006000000000000000000000000000000000000;
defparam promx9_inst_4.INIT_RAM_3A = 288'h000000000000000000000000000000000000800000000002000000000000000000000006;
defparam promx9_inst_4.INIT_RAM_3B = 288'h800000000002000000000000000000000006800000000002000000000000000000000006;
defparam promx9_inst_4.INIT_RAM_3C = 288'h800000000002000000000000000000000006800000000002000000000000000000000006;
defparam promx9_inst_4.INIT_RAM_3D = 288'h000000000778018020003008000600018000800000000002000000000000000000000006;
defparam promx9_inst_4.INIT_RAM_3E = 288'h000000000800000000002000000000000006800000000002000000000000000000000006;
defparam promx9_inst_4.INIT_RAM_3F = 288'h800000000002000000000000000000000006000000000000000000000000000000000000;

pROMX9 promx9_inst_5 (
    .DO({promx9_inst_5_dout_w[26:0],promx9_inst_5_dout[26:18]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_5.READ_MODE = 1'b0;
defparam promx9_inst_5.BIT_WIDTH = 9;
defparam promx9_inst_5.RESET_MODE = "SYNC";
defparam promx9_inst_5.INIT_RAM_00 = 288'h000000000800000AA5000018000600000000000000000800140AA00000000C0080000000;
defparam promx9_inst_5.INIT_RAM_01 = 288'h000311C00470011C0046800000000000000000000000000400000050000000030000C000;
defparam promx9_inst_5.INIT_RAM_02 = 288'h00000000000000000000000DE0000000000000000000000000000000000DE00000000000;
defparam promx9_inst_5.INIT_RAM_03 = 288'h000000000000000000000000000001BC0000000000000000000000000000000000000000;
defparam promx9_inst_5.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_5.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_5.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_5.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_5.INIT_RAM_08 = 288'h00000000000000000000000000F00180000000000000000000000000000000000000000F;
defparam promx9_inst_5.INIT_RAM_09 = 288'h00000000000000000000000000007800C000000000000000001E00300000000000000000;
defparam promx9_inst_5.INIT_RAM_0A = 288'h000000000000001E00300000000000000000000000000000001E00300000000000000000;
defparam promx9_inst_5.INIT_RAM_0B = 288'h000000000000000000F00000000000000000000000000000000000378000000000000000;
defparam promx9_inst_5.INIT_RAM_0C = 288'h000000000000000000800000000000000000000000000000000000800000000000000000;
defparam promx9_inst_5.INIT_RAM_0D = 288'h000000000000000000800000000000000000000000000000000000800000000000000000;
defparam promx9_inst_5.INIT_RAM_0E = 288'h000000000000000000800000000000000000000000000000000000E00000000000000000;
defparam promx9_inst_5.INIT_RAM_0F = 288'h00000000000000000090000000000000000000000000C02A38008E00238008D000000000;
defparam promx9_inst_5.INIT_RAM_10 = 288'h00000000000000000000400000000000000B00000000000000000000480000000000000B;
defparam promx9_inst_5.INIT_RAM_11 = 288'h00000000000000000000400000000000000B00000000000000000000480000000000000B;
defparam promx9_inst_5.INIT_RAM_12 = 288'h00000000000000000000400000000000000B00000000000000000000480000000000000B;
defparam promx9_inst_5.INIT_RAM_13 = 288'h00000000000000000000000000000000000000000000000000000000480000000000000B;
defparam promx9_inst_5.INIT_RAM_14 = 288'h00000000000000000000480000000000000B00000000000000000000480000000000000B;
defparam promx9_inst_5.INIT_RAM_15 = 288'h00000000000000000000480000000000000B00000000000000000000480000000000000B;
defparam promx9_inst_5.INIT_RAM_16 = 288'h00000000080000000500280000005A340000000000000000000000000000000000000000;
defparam promx9_inst_5.INIT_RAM_17 = 288'h000000000000000000000001E0000000000000000000000000000000780000000000000B;
defparam promx9_inst_5.INIT_RAM_18 = 288'h000000000000000000004000000000000001000000000000000000004800000000000001;
defparam promx9_inst_5.INIT_RAM_19 = 288'h000000000000000000004000000000000001000000000000000000004800000000000001;
defparam promx9_inst_5.INIT_RAM_1A = 288'h000000000000000000004000000000000001000000000000000000004800000000000001;
defparam promx9_inst_5.INIT_RAM_1B = 288'h000000100000000080001800000000000002000000000000000000004800000000000001;
defparam promx9_inst_5.INIT_RAM_1C = 288'h000000000000000000004800000000000001000000000000000000004800000000000001;
defparam promx9_inst_5.INIT_RAM_1D = 288'h000000000000000000004800000000000001000000000000000000004800000000000001;
defparam promx9_inst_5.INIT_RAM_1E = 288'h000000000800000000500011A00000000002000000000000000000000000100000014002;
defparam promx9_inst_5.INIT_RAM_1F = 288'h000000100000000080001800000000000002000000000000000000007800000000000001;
defparam promx9_inst_5.INIT_RAM_20 = 288'h000000000000000000000020000000000003000000000000000000000024000000000003;
defparam promx9_inst_5.INIT_RAM_21 = 288'h000000000000000000000020000000000003000000000000000000000024000000000003;
defparam promx9_inst_5.INIT_RAM_22 = 288'h000000000000000000000020000000000003000000000000000000000024000000000003;
defparam promx9_inst_5.INIT_RAM_23 = 288'h000020000000010000300000000000000004000000000000000000000024000000000003;
defparam promx9_inst_5.INIT_RAM_24 = 288'h000000000000000000000024000000000003000000000000000000000024000000000003;
defparam promx9_inst_5.INIT_RAM_25 = 288'h000000000000000000000024000000000003000000000000000000000024000000000003;
defparam promx9_inst_5.INIT_RAM_26 = 288'h0000001000000000A0002340000000000004000000000000000000000020000002800004;
defparam promx9_inst_5.INIT_RAM_27 = 288'h00002000000001000030000000000000000400000000000000000000003C000000000003;
defparam promx9_inst_5.INIT_RAM_28 = 288'h000000000000020000000000000000000007000000000000024000000000000000000007;
defparam promx9_inst_5.INIT_RAM_29 = 288'h000000000000020000000000000000000007000000000000024000000000000000000007;
defparam promx9_inst_5.INIT_RAM_2A = 288'h000000000000020000000000000000000007000000000000024000000000000000000007;
defparam promx9_inst_5.INIT_RAM_2B = 288'h80000000040000C000000000000000000008000000000000024000000000000000000007;
defparam promx9_inst_5.INIT_RAM_2C = 288'h000000000000024000000000000000000007000000000000024000000000000000000007;
defparam promx9_inst_5.INIT_RAM_2D = 288'h000000000000024000000000000000000007000000000000024000000000000000000007;
defparam promx9_inst_5.INIT_RAM_2E = 288'h00400000000280008D0000000000000000080000000000000000008000000A0000000008;
defparam promx9_inst_5.INIT_RAM_2F = 288'h80000000040000C00000000000000000000800000000000003C000000000000000000007;
defparam promx9_inst_5.INIT_RAM_30 = 288'h000000000000000000000020000000000009000000000000000000000024000000000009;
defparam promx9_inst_5.INIT_RAM_31 = 288'h000000000000000000000020000000000009000000000000000000000024000000000009;
defparam promx9_inst_5.INIT_RAM_32 = 288'h000000000000000000000020000000000009000000000000000000000024000000000009;
defparam promx9_inst_5.INIT_RAM_33 = 288'h00002000000001000030000000000000000A000000000000000000000024000000000009;
defparam promx9_inst_5.INIT_RAM_34 = 288'h000000000000000000000024000000000009000000000000000000000024000000000009;
defparam promx9_inst_5.INIT_RAM_35 = 288'h000000000000000000000024000000000009000000000000000000000024000000000009;
defparam promx9_inst_5.INIT_RAM_36 = 288'h0000001000000000A000234000000000000A00000000000000000000002000000280000A;
defparam promx9_inst_5.INIT_RAM_37 = 288'h00002000000001000030000000000000000A00000000000000000000003C000000000009;
defparam promx9_inst_5.INIT_RAM_38 = 288'h000000000000000000800000000000000006000000000000000000900000000000000006;
defparam promx9_inst_5.INIT_RAM_39 = 288'h000000000000000000800000000000000006000000000000000000900000000000000006;
defparam promx9_inst_5.INIT_RAM_3A = 288'h000000000000000000800000000000000006000000000000000000900000000000000006;
defparam promx9_inst_5.INIT_RAM_3B = 288'h80000000040000C000000000000000000000000000000000000000900000000000000006;
defparam promx9_inst_5.INIT_RAM_3C = 288'h000000000000000000900000000000000006000000000000000000900000000000000006;
defparam promx9_inst_5.INIT_RAM_3D = 288'h000000000000000000900000000000000006000000000000000000900000000000000006;
defparam promx9_inst_5.INIT_RAM_3E = 288'h00400000000280008D0000000000000000000000000000000000008000000A0000000000;
defparam promx9_inst_5.INIT_RAM_3F = 288'h80000000040000C000000000000000000000000000000000000000F00000000000000006;

pROMX9 promx9_inst_6 (
    .DO({promx9_inst_6_dout_w[26:0],promx9_inst_6_dout[35:27]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_6.READ_MODE = 1'b0;
defparam promx9_inst_6.BIT_WIDTH = 9;
defparam promx9_inst_6.RESET_MODE = "SYNC";
defparam promx9_inst_6.INIT_RAM_00 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_01 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_02 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_03 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_04 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_05 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_06 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_07 = 288'h0000000000000000023A00000020400000040000000000000000023A0000002040000004;
defparam promx9_inst_6.INIT_RAM_08 = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_09 = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_0A = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_0B = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_0C = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_0D = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_0E = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_0F = 288'h000000000004000002040000000000000004000000000004000002040000000000000004;
defparam promx9_inst_6.INIT_RAM_10 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_11 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_12 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_13 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_14 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_15 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_16 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_17 = 288'h000000000000000000000000474000000008000000000000000000000000474000000008;
defparam promx9_inst_6.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000004000064298000000000000008;
defparam promx9_inst_6.INIT_RAM_19 = 288'h000000000004000004298000000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000004000004290000000000000008;
defparam promx9_inst_6.INIT_RAM_1B = 288'h000000000004000004290000000000000008000000000004000004290000000000000008;
defparam promx9_inst_6.INIT_RAM_1C = 288'h000000000004000004290000000000000008000000000004000004290000000000000008;
defparam promx9_inst_6.INIT_RAM_1D = 288'h00000000000000000000000000000400C882000000000004000064290000000000000008;
defparam promx9_inst_6.INIT_RAM_1E = 288'h0000000000000000000000000A4290000008000000000004000064290000000000000008;
defparam promx9_inst_6.INIT_RAM_1F = 288'h000000000004000004510000000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000001902600000000000000000008;
defparam promx9_inst_6.INIT_RAM_21 = 288'h000000000000102600000000000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000102400000000000000000008;
defparam promx9_inst_6.INIT_RAM_23 = 288'h000000000000102400000000000000000008000000000000102400000000000000000008;
defparam promx9_inst_6.INIT_RAM_24 = 288'h000000000000102400000000000000000008000000000000102400000000000000000008;
defparam promx9_inst_6.INIT_RAM_25 = 288'h00000000000000000000000010041400C882000000000001902400000000000000000008;
defparam promx9_inst_6.INIT_RAM_26 = 288'h000000000002902400000000000000000008000000000001902400000000000000000008;
defparam promx9_inst_6.INIT_RAM_27 = 288'h000000000000114400000000000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000001912600000000000000000008;
defparam promx9_inst_6.INIT_RAM_29 = 288'h000000000000112600000000000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000112400000000000000000008;
defparam promx9_inst_6.INIT_RAM_2B = 288'h000000000000112400000000000000000008000000000000112400000000000000000008;
defparam promx9_inst_6.INIT_RAM_2C = 288'h000000000000112400000000000000000008000000000000112400000000000000000008;
defparam promx9_inst_6.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000001912400000000000000000008;
defparam promx9_inst_6.INIT_RAM_2E = 288'h000000000002912400000000000000000008000000000001912400000000000000000008;
defparam promx9_inst_6.INIT_RAM_2F = 288'h000000000000114400000000000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_30 = 288'h0000000000000000000000000000000000000000000000000200003214C0000000000008;
defparam promx9_inst_6.INIT_RAM_31 = 288'h0000000000000200000214C0000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000020000021480000000000008;
defparam promx9_inst_6.INIT_RAM_33 = 288'h000000000000020000021480000000000008000000000000020000021480000000000008;
defparam promx9_inst_6.INIT_RAM_34 = 288'h000000000000020000021480000000000008000000000000020000021480000000000008;
defparam promx9_inst_6.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000020000321480000000000008;
defparam promx9_inst_6.INIT_RAM_36 = 288'h000000000000000000000000000521480008000000000000020000321480000000000008;
defparam promx9_inst_6.INIT_RAM_37 = 288'h000000000000020000022880000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_38 = 288'h00000000000000000000000000000000000000000000080000C853000000000000000008;
defparam promx9_inst_6.INIT_RAM_39 = 288'h000000000800000853000000000000000008000000000000000000000000000000000000;
defparam promx9_inst_6.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000800000852000000000000000008;
defparam promx9_inst_6.INIT_RAM_3B = 288'h000000000800000852000000000000000008000000000800000852000000000000000008;
defparam promx9_inst_6.INIT_RAM_3C = 288'h000000000800000852000000000000000008000000000800000852000000000000000008;
defparam promx9_inst_6.INIT_RAM_3D = 288'h00000000041008008201001040200208000000000000080000C852000000000000000008;
defparam promx9_inst_6.INIT_RAM_3E = 288'h00000000000000000000001485200000000800000000080000C852000000000000000008;
defparam promx9_inst_6.INIT_RAM_3F = 288'h0000000008000008A2000000000000000008000000000000000000000000000000000000;

pROMX9 promx9_inst_7 (
    .DO({promx9_inst_7_dout_w[26:0],promx9_inst_7_dout[35:27]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_7.READ_MODE = 1'b0;
defparam promx9_inst_7.BIT_WIDTH = 9;
defparam promx9_inst_7.RESET_MODE = "SYNC";
defparam promx9_inst_7.INIT_RAM_00 = 288'h000000000000000000010000082001900082000000000000000000010010400410000064;
defparam promx9_inst_7.INIT_RAM_01 = 288'h00000002200048009200000000000000007200000000000000000000008000000000C842;
defparam promx9_inst_7.INIT_RAM_02 = 288'h000000000000000000000000094010001000000000000000000000000000002000200008;
defparam promx9_inst_7.INIT_RAM_03 = 288'h000000000000000000000000000000000408000000000000000000000000000000000000;
defparam promx9_inst_7.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_7.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_7.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_7.INIT_RAM_07 = 288'h000000000000000000000000000000000008000000000000000000000000000000000008;
defparam promx9_inst_7.INIT_RAM_08 = 288'h000000000000000000000000000000000408000000000000000000000000000000000008;
defparam promx9_inst_7.INIT_RAM_09 = 288'h000000000000000000000000000000000092000000000000000000000080000000200008;
defparam promx9_inst_7.INIT_RAM_0A = 288'h000000000000000000002500400040001000000000000000000000002500400000001000;
defparam promx9_inst_7.INIT_RAM_0B = 288'h000000000000000000000102400000000008000000000000000000002500400040001000;
defparam promx9_inst_7.INIT_RAM_0C = 288'h000000000000000000000100400000000008000000000000000000000100400000000008;
defparam promx9_inst_7.INIT_RAM_0D = 288'h000000000000000000000100400000000008000000000000000000000100400000000008;
defparam promx9_inst_7.INIT_RAM_0E = 288'h000000000000000000000100400000000008000000000000000000000114600000000008;
defparam promx9_inst_7.INIT_RAM_0F = 288'h000000000000000000000112400000000008000000000000004400090012400000000072;
defparam promx9_inst_7.INIT_RAM_10 = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_11 = 288'h00000000000000000000000A89200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_12 = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000852000000008;
defparam promx9_inst_7.INIT_RAM_14 = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_15 = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_16 = 288'h00000000000000000000000047400000E46C000000000000000000000000000000000000;
defparam promx9_inst_7.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000852000000008;
defparam promx9_inst_7.INIT_RAM_18 = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_19 = 288'h00000000000000000000000A89200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_1A = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_1B = 288'h00000000000002000009000A400000000008000000000000000000000000852000000008;
defparam promx9_inst_7.INIT_RAM_1C = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_1D = 288'h00000000000000000000000A81200000000800000000000000000000000A812000000008;
defparam promx9_inst_7.INIT_RAM_1E = 288'h000000000000000000000C80072000000008000000000000000000000000000000000008;
defparam promx9_inst_7.INIT_RAM_1F = 288'h00000000000002000049000A400000000008000000000000000000000000852000000008;
defparam promx9_inst_7.INIT_RAM_20 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_21 = 288'h000000000000000000000000054490000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_22 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_23 = 288'h000000000004000012000C80000000000008000000000000000000000000004290000008;
defparam promx9_inst_7.INIT_RAM_24 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_25 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_26 = 288'h00000000000000000019000E400000000008000000000000000000000000000000006408;
defparam promx9_inst_7.INIT_RAM_27 = 288'h000000000004000092000C80000000000008000000000000000000000000004290000008;
defparam promx9_inst_7.INIT_RAM_28 = 288'h000000000000000054090000000000000008000000000000000054090000000000000008;
defparam promx9_inst_7.INIT_RAM_29 = 288'h000000000000000054490000000000000008000000000000000054090000000000000008;
defparam promx9_inst_7.INIT_RAM_2A = 288'h000000000000000054090000000000000008000000000000000054090000000000000008;
defparam promx9_inst_7.INIT_RAM_2B = 288'h000000100000480032000000000000000008000000000000000004290000000000000008;
defparam promx9_inst_7.INIT_RAM_2C = 288'h000000000000000054090000000000000008000000000000000054090000000000000008;
defparam promx9_inst_7.INIT_RAM_2D = 288'h000000000000000054090000000000000008000000000000000054090000000000000008;
defparam promx9_inst_7.INIT_RAM_2E = 288'h000000000000006400390000000000000008000000000000000000000000000190000008;
defparam promx9_inst_7.INIT_RAM_2F = 288'h000000100002480032000000000000000008000000000000000004290000000000000008;
defparam promx9_inst_7.INIT_RAM_30 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_31 = 288'h000000000000000000000000054490000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_32 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_33 = 288'h000000000004000012000C80000000000008000000000000000000000000004290000008;
defparam promx9_inst_7.INIT_RAM_34 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_35 = 288'h000000000000000000000000054090000008000000000000000000000000054090000008;
defparam promx9_inst_7.INIT_RAM_36 = 288'h00000000000000000019000E400000000008000000000000000000000000000000006408;
defparam promx9_inst_7.INIT_RAM_37 = 288'h000000000004000092000C80000000000008000000000000000000000000004290000008;
defparam promx9_inst_7.INIT_RAM_38 = 288'h000000000000000000001502400000000008000000000000000000001502400000000008;
defparam promx9_inst_7.INIT_RAM_39 = 288'h000000000000000000001512400000000008000000000000000000001502400000000008;
defparam promx9_inst_7.INIT_RAM_3A = 288'h000000000000000000001502400000000008000000000000000000001502400000000008;
defparam promx9_inst_7.INIT_RAM_3B = 288'h00000010000048009200000000000000000800000000000000000000010A400000000008;
defparam promx9_inst_7.INIT_RAM_3C = 288'h000000000000000000001502400000000008000000000000000000001502400000000008;
defparam promx9_inst_7.INIT_RAM_3D = 288'h000000000000000000001502400000000008000000000000000000001502400000000008;
defparam promx9_inst_7.INIT_RAM_3E = 288'h000000000000012400390000000000000008000000000000000000000000000490000008;
defparam promx9_inst_7.INIT_RAM_3F = 288'h00000010000248009200000000000000000800000000000000000000010A400000000008;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[27:0],dout[39:36]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_8.READ_MODE = 1'b0;
defparam prom_inst_8.BIT_WIDTH = 4;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_12 = 256'h0000000000020000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_20 = 256'h0100000000000000000000000020000000000000020000000000000002000000;
defparam prom_inst_8.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000200;
defparam prom_inst_8.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_23 = 256'h0000000000000000000000000000000400000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_24 = 256'h0000000000000000000000000000020000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_25 = 256'h0000000000000000000000000000200000000000000020000000000000000000;
defparam prom_inst_8.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(promx9_inst_0_dout[0]),
  .I1(promx9_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(promx9_inst_0_dout[1]),
  .I1(promx9_inst_1_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_2 (
  .O(dout[2]),
  .I0(promx9_inst_0_dout[2]),
  .I1(promx9_inst_1_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(dout[3]),
  .I0(promx9_inst_0_dout[3]),
  .I1(promx9_inst_1_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_4 (
  .O(dout[4]),
  .I0(promx9_inst_0_dout[4]),
  .I1(promx9_inst_1_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[5]),
  .I0(promx9_inst_0_dout[5]),
  .I1(promx9_inst_1_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_6 (
  .O(dout[6]),
  .I0(promx9_inst_0_dout[6]),
  .I1(promx9_inst_1_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_7 (
  .O(dout[7]),
  .I0(promx9_inst_0_dout[7]),
  .I1(promx9_inst_1_dout[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[8]),
  .I0(promx9_inst_0_dout[8]),
  .I1(promx9_inst_1_dout[8]),
  .S0(dff_q_0)
);
MUX2 mux_inst_9 (
  .O(dout[9]),
  .I0(promx9_inst_2_dout[9]),
  .I1(promx9_inst_3_dout[9]),
  .S0(dff_q_0)
);
MUX2 mux_inst_10 (
  .O(dout[10]),
  .I0(promx9_inst_2_dout[10]),
  .I1(promx9_inst_3_dout[10]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[11]),
  .I0(promx9_inst_2_dout[11]),
  .I1(promx9_inst_3_dout[11]),
  .S0(dff_q_0)
);
MUX2 mux_inst_12 (
  .O(dout[12]),
  .I0(promx9_inst_2_dout[12]),
  .I1(promx9_inst_3_dout[12]),
  .S0(dff_q_0)
);
MUX2 mux_inst_13 (
  .O(dout[13]),
  .I0(promx9_inst_2_dout[13]),
  .I1(promx9_inst_3_dout[13]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[14]),
  .I0(promx9_inst_2_dout[14]),
  .I1(promx9_inst_3_dout[14]),
  .S0(dff_q_0)
);
MUX2 mux_inst_15 (
  .O(dout[15]),
  .I0(promx9_inst_2_dout[15]),
  .I1(promx9_inst_3_dout[15]),
  .S0(dff_q_0)
);
MUX2 mux_inst_16 (
  .O(dout[16]),
  .I0(promx9_inst_2_dout[16]),
  .I1(promx9_inst_3_dout[16]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[17]),
  .I0(promx9_inst_2_dout[17]),
  .I1(promx9_inst_3_dout[17]),
  .S0(dff_q_0)
);
MUX2 mux_inst_18 (
  .O(dout[18]),
  .I0(promx9_inst_4_dout[18]),
  .I1(promx9_inst_5_dout[18]),
  .S0(dff_q_0)
);
MUX2 mux_inst_19 (
  .O(dout[19]),
  .I0(promx9_inst_4_dout[19]),
  .I1(promx9_inst_5_dout[19]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(dout[20]),
  .I0(promx9_inst_4_dout[20]),
  .I1(promx9_inst_5_dout[20]),
  .S0(dff_q_0)
);
MUX2 mux_inst_21 (
  .O(dout[21]),
  .I0(promx9_inst_4_dout[21]),
  .I1(promx9_inst_5_dout[21]),
  .S0(dff_q_0)
);
MUX2 mux_inst_22 (
  .O(dout[22]),
  .I0(promx9_inst_4_dout[22]),
  .I1(promx9_inst_5_dout[22]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(dout[23]),
  .I0(promx9_inst_4_dout[23]),
  .I1(promx9_inst_5_dout[23]),
  .S0(dff_q_0)
);
MUX2 mux_inst_24 (
  .O(dout[24]),
  .I0(promx9_inst_4_dout[24]),
  .I1(promx9_inst_5_dout[24]),
  .S0(dff_q_0)
);
MUX2 mux_inst_25 (
  .O(dout[25]),
  .I0(promx9_inst_4_dout[25]),
  .I1(promx9_inst_5_dout[25]),
  .S0(dff_q_0)
);
MUX2 mux_inst_26 (
  .O(dout[26]),
  .I0(promx9_inst_4_dout[26]),
  .I1(promx9_inst_5_dout[26]),
  .S0(dff_q_0)
);
MUX2 mux_inst_27 (
  .O(dout[27]),
  .I0(promx9_inst_6_dout[27]),
  .I1(promx9_inst_7_dout[27]),
  .S0(dff_q_0)
);
MUX2 mux_inst_28 (
  .O(dout[28]),
  .I0(promx9_inst_6_dout[28]),
  .I1(promx9_inst_7_dout[28]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(dout[29]),
  .I0(promx9_inst_6_dout[29]),
  .I1(promx9_inst_7_dout[29]),
  .S0(dff_q_0)
);
MUX2 mux_inst_30 (
  .O(dout[30]),
  .I0(promx9_inst_6_dout[30]),
  .I1(promx9_inst_7_dout[30]),
  .S0(dff_q_0)
);
MUX2 mux_inst_31 (
  .O(dout[31]),
  .I0(promx9_inst_6_dout[31]),
  .I1(promx9_inst_7_dout[31]),
  .S0(dff_q_0)
);
MUX2 mux_inst_32 (
  .O(dout[32]),
  .I0(promx9_inst_6_dout[32]),
  .I1(promx9_inst_7_dout[32]),
  .S0(dff_q_0)
);
MUX2 mux_inst_33 (
  .O(dout[33]),
  .I0(promx9_inst_6_dout[33]),
  .I1(promx9_inst_7_dout[33]),
  .S0(dff_q_0)
);
MUX2 mux_inst_34 (
  .O(dout[34]),
  .I0(promx9_inst_6_dout[34]),
  .I1(promx9_inst_7_dout[34]),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(dout[35]),
  .I0(promx9_inst_6_dout[35]),
  .I1(promx9_inst_7_dout[35]),
  .S0(dff_q_0)
);
endmodule //Gowin_pROM_uc
