
library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_apple2 is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM_apple2;

architecture Behavioral of Gowin_pROM_apple2 is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"80108C416F80258C0085C82F7E10A237800040D0BF7570A2A5E5EA881A1A2262",
            INIT_RAM_02 => X"0092864EF256D4188B6F7E14091088F6080CC0002B3599C0B2024B6441005120",
            INIT_RAM_03 => X"683338CEA246C570385C241EB028C8C8261A440209A69900C34266D181E80802",
            INIT_RAM_04 => X"494BD404D6BAA67E175CC652402040CE302D4802129906890260990B249A0008",
            INIT_RAM_05 => X"3082B2D6239820202112587996408004286A6D1EAB3D5C9C7D7A80F2121B00F4",
            INIT_RAM_06 => X"5253496068C8C4D10859189400CD0F3DCBB68801A1E7B62EDA089126241A8D01",
            INIT_RAM_07 => X"6DFF19509C000DFDFDF25A3170B94D23080A5880421604FAB3817D422904F6CC",
            INIT_RAM_08 => X"CA583402C306A2EF7AB034071501503600626C5DE91F806303DFDC60DB80F804",
            INIT_RAM_09 => X"02433858F4100DB640338CE125B6586AA44780C07926EA62E3F0A98090D1AA9E",
            INIT_RAM_0A => X"3E4BE05AC390A38B7098C0486611040082249EDA8090DFD8F89105FECE960430",
            INIT_RAM_0B => X"8C4F1595FE89BE0E5E588CBA8391D6391AD7F4EEA4FADBF618C43123233E6703",
            INIT_RAM_0C => X"0B0B4C210151441809405192BA0698F8218106028A4548B184843FAA281CA690",
            INIT_RAM_0D => X"C47000028E02C0884C008128207079522BBA25F3FC9066BB6503AD21BF112F25",
            INIT_RAM_0E => X"3B07FEF05BE00F05AC602050308392060066220020C21C9060008C25B3329247",
            INIT_RAM_0F => X"E332290E220840256F02F2C4E00410D09D921A0205C64A110C09A8A689278F0A",
            INIT_RAM_10 => X"87612D9268918DC84FF501F20EF97036344A4F7A8BD6F158402A6A4F12EBEB8D",
            INIT_RAM_11 => X"B54A29166D63272B675714F5655AB6A77C579E455B34B5CB8CEF5C98C4564488",
            INIT_RAM_12 => X"47348F593A2D91D4A6F278B4E7344DE66293466218C21E85714F9C1E038E9692",
            INIT_RAM_13 => X"680C86000C8296290AA94C1CE8F0257BBFA37C0F22526A29D32D3B2D53295F53",
            INIT_RAM_14 => X"9268DE33D674A1DCCC22A2A949E2EBEDEBFC0B00A58208892D092A20C4A25C00",
            INIT_RAM_15 => X"703A688B315F9663AF930C0021F691938512888080E299FF0B148313A12405F9",
            INIT_RAM_16 => X"994079903B7340213101260F5F1500123333314ABEFB2C5983323CB38CF7A580",
            INIT_RAM_17 => X"A56824860901B2A6469589B5DD06C9C9A61AC1461291292289860931B359D493",
            INIT_RAM_18 => X"25910A16577720B21ABE19CE2082AC333048B516591A3CA4213066205A34E010",
            INIT_RAM_19 => X"02B101254B0DAC14844E420214D92E04012DF357C06292D8244592E782812726",
            INIT_RAM_1A => X"9AD2B186630B35AD149C39C8A6D82354A33DA480C66427828763D50137FA0042",
            INIT_RAM_1B => X"393C5A4A4466764D8685969449C3441199060DEC5CC968C018C902C8680A29A3",
            INIT_RAM_1C => X"40A6AAD1A1D8A8D54296A4068784A4CE74C920105B2653B39A2A944914784282",
            INIT_RAM_1D => X"306E2028532444FAEE28BBF7765A260100A5432528D3ED6FEE4B43794000418F",
            INIT_RAM_1E => X"44808900A9D880A44BCA4C9C2B01D9333362212D7AB2CB252641965C30815306",
            INIT_RAM_1F => X"44292C4050345B1114A2213C664098C5B10D76DA1677C0FE83000B20C890B188",
            INIT_RAM_20 => X"128F6342F6DB3AF0D3A569333033563762F0C9E6181AC12508BD46CF11492904",
            INIT_RAM_21 => X"B3260363834BE4E40956681904A73634D942CCEB0853F5750B464196610679C8",
            INIT_RAM_22 => X"62615E02D53122000DF38CED04057256090D0960790EF874E7A8A5427849D90C",
            INIT_RAM_23 => X"3352643811019084444464A596674A5E0332699405E93143B16C822655301402",
            INIT_RAM_24 => X"084F4A88932E27E6D6127F6993338661A0E0676423680A40FAE282164888F499",
            INIT_RAM_25 => X"80F06820CCCC01C1330258B40585C5524F5771E850AFE6588120514853612A17",
            INIT_RAM_26 => X"265B10046C101E4181778808035E348442809C042808D887A608079510444299",
            INIT_RAM_27 => X"AB4AC081C20C383581BD77411A849142265891964C3C09904809492A50140828",
            INIT_RAM_28 => X"4241828208408081DFDDFDD744411FD82234AFEAFEA74520A08004EF4BBD2BA2",
            INIT_RAM_29 => X"D5695A4808857F57F442199C671DD44B4A4B93AC4CBD7E88A02D4843B3080454",
            INIT_RAM_2A => X"923D7D4408020AFEAFE008861A280280C21E619281C054810C8169C5A11ADE95",
            INIT_RAM_2B => X"D08E626BA51A95A14124259D69AC666D022C45208B2872E9CA72210406955A56",
            INIT_RAM_2C => X"042865D6B9892288170A850E6A090111899C8C65647480DD5FA44838CA280381",
            INIT_RAM_2D => X"3CA0DC0016E75B9613219A129672E9091209212FF4C0AA52C0E92099D24E6529",
            INIT_RAM_2E => X"38C2DE03C9D30D871A5054E01621DE0E864A0804D595AEC92FF240D22701D4C9",
            INIT_RAM_2F => X"C03D0710D753693A6231108430D63C605F0F1CDE306C11165DCD6D29E325C611",
            INIT_RAM_30 => X"840D61E3071F4261B41176C44463BBFB662139D008551E0CBA189043B323866A",
            INIT_RAM_31 => X"0024040804C8C665630B01033382E2EC4895FAF281343B5D549CA23129130063",
            INIT_RAM_32 => X"EBEBC126B8F5187D1F47D98BFA27D9A3499808C3480004048008408003350991",
            INIT_RAM_33 => X"4354B50442585E716594AF3B631910442FC0138B5C4003AE0054A2F57D913EFA",
            INIT_RAM_34 => X"985158E406C07F505474E4BCE00724E8996058C5550516ACD0DF121945423E01",
            INIT_RAM_35 => X"6330D1B5CD0BCDDA8406F548C82ABBAA4AFCA17124AFD78F10EA845454842CE6",
            INIT_RAM_36 => X"F3090018500211114C1801C56E029A0D086646C101801C16E429A0D086646C10",
            INIT_RAM_37 => X"90266805CA0E4423F2D8884CC4F11984630B2CD2168F452908F5082124481A4A",
            INIT_RAM_38 => X"05396814A5101C08F0C03482A62219218050507C94716E005A8960C0805554C8",
            INIT_RAM_39 => X"7AF5183CEED6FDF804AC7198646664606060644094B0668844159135F7022836",
            INIT_RAM_3A => X"211DE39B5E020ED9EB19CD2091DAD7F03A44A58301328CCF0000000000000000",
            INIT_RAM_3B => X"234442102651C5B82320263B10615015035FA1F01FB0AA19964A80206BF9A2EA",
            INIT_RAM_3C => X"31EF6C0899856683D6018C840C81CF1EEA188F94324840A030C3141E34709131",
            INIT_RAM_3D => X"011208BB01B388008E65BEEEC90AC19093C96E66481923124B9B24A89024A666",
            INIT_RAM_3E => X"602484942711B0210C90218268290A22458B270290DC7398C15054567C40BC88",
            INIT_RAM_3F => X"8FD7F895CB19046E72CA5013F3100B10A236DB0960448C8CEF6772E23257460E"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"54804422557080B50C0080AA0002A1210D2012C28A0300046101119004100606",
            INIT_RAM_02 => X"34830A8A00008084920A21920080045D6028816120AD02A20100120A08249300",
            INIT_RAM_03 => X"41020808C0A08640288413311DC08410041EE6029114110189104411136CA016",
            INIT_RAM_04 => X"15A2C484485A062E4009B0202761352200091840012621401000214000000300",
            INIT_RAM_05 => X"48150A4204A085050400C851021A0500800081000A2088502800151001F04080",
            INIT_RAM_06 => X"54480010B448AC2084C324331B1408A10024463681142400915F608108088420",
            INIT_RAM_07 => X"6150459CD92960D491720C095D0120003A62418346954CD6AE28352A14E41851",
            INIT_RAM_08 => X"821365818624124A521261A21511510C24C0240829088001D882A920804884A0",
            INIT_RAM_09 => X"B2266E93A5308804220AD83001084C34C6A6C402500C08485A500148A588A094",
            INIT_RAM_0A => X"1842C548C3181940280840000008248866AB3491B57094B611871D8C44024291",
            INIT_RAM_0B => X"604322F521092C0E5E3589BA92891524C4909A4124908D134000102112284403",
            INIT_RAM_0C => X"404808E0801050A0608700104A064285682490541002011041B4B446F99329D2",
            INIT_RAM_0D => X"1214442002900DD00118400AAD1A525211010881000A45204890202C0A890425",
            INIT_RAM_0E => X"B4208C6E150099091A200402022011405154112808088082540844012A802232",
            INIT_RAM_0F => X"E02804C18104FDCAE294B02265128D4410A94248084414C710003154000B0DC3",
            INIT_RAM_10 => X"83B06200807A9FF9A992FEEE5B8EE776BA2F4D14802BFEA7FFAE7EABA80BAA09",
            INIT_RAM_11 => X"D1642F253147534521D4E37B5AD805A28BB8A094DA5B0EAD44866514A436DD30",
            INIT_RAM_12 => X"821A5A86211E8A04C9863B610200C6E22C45E22100A45C5644978CEE0F7B2E75",
            INIT_RAM_13 => X"0C585402B155C810843A94495230CC894854002CC47CCD3227341B03F3354402",
            INIT_RAM_14 => X"14508A88483028A08895C13A284950090450684D702F2114E12D18226D211102",
            INIT_RAM_15 => X"1A12A9428209004582080472A28000220A028D028A80C2A561D2DAE14628028A",
            INIT_RAM_16 => X"0C10133020280A00016800420A081468828228C411524053220220A61848B05E",
            INIT_RAM_17 => X"08001410300C053214A14AAAA4A01000B07498025090A96A0301CD08E6103592",
            INIT_RAM_18 => X"AA0052A0A802410400144100AB80A0288180291A1040092B000400B0184CA64C",
            INIT_RAM_19 => X"412040A5208124050831A15980404288B7184000ACC242253240203424995004",
            INIT_RAM_1A => X"86C01102400A00002000208182008A14130000D0120A11B0601420FC08295220",
            INIT_RAM_1B => X"208C60246450236D2529884E046298241110010A084909519AD854D910216022",
            INIT_RAM_1C => X"40498788B150A491080421D2C1348088244B4842D2002054008000CD07211213",
            INIT_RAM_1D => X"00A259DAD0148B4A2A1000095441308ACAC501200B380280A0C3688608108923",
            INIT_RAM_1E => X"8134206510C81220005A54A8080298015004050015009054A2482406270E8884",
            INIT_RAM_1F => X"5AC8214853A6D8ACDD02E952008C0B221382AA10101021421B24408658852900",
            INIT_RAM_20 => X"0008C204A492148081804A822054B40400A09114126050A06242220288430000",
            INIT_RAM_21 => X"2A0801C27A921860B0C4408852E264AA110466504A1008029020802235880240",
            INIT_RAM_22 => X"669604121304AD1710214808E1EA0D692642055540905221541360191A4401D3",
            INIT_RAM_23 => X"02545B8B4231084888880125224084062204D522C9455825800821160DA248C0",
            INIT_RAM_24 => X"90C081131CA29292041D9522E46C833100930501024D8C09440B2D1C5061202A",
            INIT_RAM_25 => X"0E00112C9880A12802241020800838191A0A842C7D48BB8C88AA265085280FA8",
            INIT_RAM_26 => X"420220828904001009110272684521127504089011108385440B3515109884A0",
            INIT_RAM_27 => X"29220060A8810774810AA968041C92E07400180006826C832048008723C8AA24",
            INIT_RAM_28 => X"202008A2052EE6648208AAAA8AFCC142F54155400048001577EC150291200508",
            INIT_RAM_29 => X"AA50845295FAAA00002AC2100000A3290062818B160040ACC0210DD39F002FAB",
            INIT_RAM_2A => X"14802A9387F19554000ABD6040800A8A19C034A4D8C04EDA1C10529400020122",
            INIT_RAM_2B => X"A42254012050200A08018840D31615814A6090F120D085529082F48641229421",
            INIT_RAM_2C => X"19800A8D5980046904723850AB108031044402A04615300A00128C0055900860",
            INIT_RAM_2D => X"AA20A8D4295A3040821522AD2D441D064CAC558890106904840C21E61077AD40",
            INIT_RAM_2E => X"66517FB162A8A888105895631048DF0E86828E0001005551C00C0B840444B094",
            INIT_RAM_2F => X"DB2D8B0A008C9D4AAC03A2061A00851C11A11654844689888021016835A05402",
            INIT_RAM_30 => X"19CAC07706ABD262842C5024B03EA5616D81EF1312A216391204982545058342",
            INIT_RAM_31 => X"120C499B0642002B626E418910004042006806A07A89208830407F7008A8C83F",
            INIT_RAM_32 => X"10546E1542009480A0008C8050280C86735305B347060018083041089040000A",
            INIT_RAM_33 => X"228029001098442A49A2426A411246831432D9000B332005A6BD3700A2C95100",
            INIT_RAM_34 => X"748894817085A8AE0A005910000010444028024A2000812841AAFFF2B80CAB8A",
            INIT_RAM_35 => X"18428E4ABAF6B4001C08000AA4504010100A3AA210008128810032A20A00E044",
            INIT_RAM_36 => X"2A8689842120204264AECE1110000D52D22C2DBF6AECE1110400D52D22C2DBF6",
            INIT_RAM_37 => X"B6710600C00420284200810A102AA2008212480480B89A3A53888E1913124250",
            INIT_RAM_38 => X"2A04011892A214384D42CA005C44A0AD78920F282BA8452008A8002400A8A289",
            INIT_RAM_39 => X"4280030E2E882A6A008382342828282820202C0021A083540AA2514402B2E044",
            INIT_RAM_3A => X"40A00C0C01000848104BA330D18B50D836084DA265248160463F5C8EB8800036",
            INIT_RAM_3B => X"08100000140CA014020911434041501500432280451010908010001821F500E8",
            INIT_RAM_3C => X"9128A410C24A246623B400050541209823226840300840AA0820000109010A81",
            INIT_RAM_3D => X"D000551078015742401511400092004C801A890268809C424A10450190E0A550",
            INIT_RAM_3E => X"412092890409124B2D10640051C130AA18A82901000280042210852908324559",
            INIT_RAM_3F => X"FEC3FE2BC6B1E00CB4511ED0283FFF18823655936830B0B00808103800030290"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0CCC6AD0CE082211A08086432D3227DEC24FED2DB912E8004482AB0D9B081479",
            INIT_RAM_02 => X"38CC84060486B00D0B765D18890C887E660A80153836A181030455004105E22A",
            INIT_RAM_03 => X"6E9190C6666643301058767FE8905CC8621E8046029A68B342422A5682978405",
            INIT_RAM_04 => X"0C63D19946307C50041804200001B4261E414C070225330688E618990C820000",
            INIT_RAM_05 => X"70A7D084A7A83021292458799440808C2842881FE8B7D4C4F53B81B8338A6CF0",
            INIT_RAM_06 => X"10492330B4704A41AAC970432047052480926440E0A4930249E57984141C8E11",
            INIT_RAM_07 => X"2E3711E0E934B1E021024C1A789124813C00008346450CF4AA21210830049284",
            INIT_RAM_08 => X"482B5181750B83B6A06A56222013012A20A35A54D2F72063991B39D8D9414C31",
            INIT_RAM_09 => X"C5325029619CCD9A0800744534B830C70C159813B13A60A00A10916C214D682D",
            INIT_RAM_0A => X"1405A122A28CA30180118B6D6243040000046D68D5356D68E9430D5A8A0D4068",
            INIT_RAM_0B => X"86668768DF82D261800E412ACDA2905FDA036FA6816816A542042A10055AA001",
            INIT_RAM_0C => X"0A0E54608C6004083C610898343AF87F49C1B248012C2011C3022AAC109A0260",
            INIT_RAM_0D => X"C66324160C08408ACCC02C306030B3C328880CE23698AB58A6098931F609AB86",
            INIT_RAM_0E => X"8D175AD4AB40968E175002C03891987070B4013580E248C242086A02A0828345",
            INIT_RAM_0F => X"DA81E1C672AC2A024C823080EA77D997C9125D9001621A07C009B15E04889204",
            INIT_RAM_10 => X"D885B57E96DFFFFDC092EFDF4A8F79189B58484040511151517EFEE10551206D",
            INIT_RAM_11 => X"A6F6878FE69EC57CB9DB5CBDAB7FF2D97477DC3570E7571E3671DC529E5C4575",
            INIT_RAM_12 => X"2BD418A0768127E9FCF6FEEB4BCADD6EAB8C6EAB6E9F816BB6B11F82C8A46DDD",
            INIT_RAM_13 => X"6B04070ADD03E8559FB3D83DBBC00478E72604092452D77FEE71B39DFBB2294D",
            INIT_RAM_14 => X"1EF8035F6D4637F5F421C13320A6CAA0BEE14E25772E815D0830121080461D20",
            INIT_RAM_15 => X"5A00EDC108001C55AB0A0660B3B3A88AA389CB8362B088E6091443E1C30975D2",
            INIT_RAM_16 => X"C9C320008169410A814550065B340030FD57D0CA3A7264400820048D1CCA254C",
            INIT_RAM_17 => X"AC62040B3508378614805FAF9D20D84810124B014AC88D2ECD258AAB404384CA",
            INIT_RAM_18 => X"FCF0BCF0D55761C60ABE7BAB44BD087F59AC023401784D61900202280B7A2728",
            INIT_RAM_19 => X"290842C52B9428002C3FF32114096C0B4C05D1346CF25074AA41B250F719EBEE",
            INIT_RAM_1A => X"535A644A1049294A3796DF40D6585B1481A52200C4261F08475575D98DE94290",
            INIT_RAM_1B => X"75F8F93F82073906A12002022A8A34AFED4645640A304500884C428819010832",
            INIT_RAM_1C => X"04BEBB858D504DEC01822000767095DD4948301519017591D88C42A1046D7257",
            INIT_RAM_1D => X"4024511A5B240DDC689A1140144910228D202A60481529CEE2216F48080004BE",
            INIT_RAM_1E => X"2048012C959CA840A49383024302E80B11152A046A92DB67084DB6483785BD80",
            INIT_RAM_1F => X"6A512542518A843015126137062E5FE2940BE4C48767D0E71384093690802A01",
            INIT_RAM_20 => X"1E366D18400002135E3C4FFDD0145421109208236E2E46C320152C86A9002879",
            INIT_RAM_21 => X"80000803C0406C054B2168392D2C10864177BAC94C90A51109024096CC0839C0",
            INIT_RAM_22 => X"93D35ED042330F8004C665E72304367B890F5705091E604D83BBC979E019DDFE",
            INIT_RAM_23 => X"B85FBE3F9EA1188000002544962D0848C0602094848AB320D125A124C88530E1",
            INIT_RAM_24 => X"100F9F111F4EFF3C937EBD49F2DF47D09860AE7187448528EEF6A66A05E3D603",
            INIT_RAM_25 => X"C450103C000F36EDF952019684D1E323DF3D126479EDD7F46B3A62109443BF3E",
            INIT_RAM_26 => X"4604A0C263900EC089231012684D692E6786F40A52904102236F2787208886F5",
            INIT_RAM_27 => X"A53A3290972D39C82175647A1E1E11E031481092A80EE98BE088008773FAB334",
            INIT_RAM_28 => X"3620755DF2CCE46FB659EFB65AF9D958F5C7FFEAABA720DD77CC11A342875B22",
            INIT_RAM_29 => X"56718D7A3F575DDF70046B18423F51101662C181062C5900805AC0940E011AAA",
            INIT_RAM_2A => X"5EDDF76CD810DFFEAAA2BD61181653CF235E040840015E4000D94949955ADF31",
            INIT_RAM_2B => X"820CC22704183031201497D45998044D8ACD8F831F2BB5CAD29BC7C11F319C63",
            INIT_RAM_2C => X"043381BAA01700454222140A45A8B87401440A811350405F3B81701B5F89888B",
            INIT_RAM_2D => X"A8D08A0539F362E21A112C0A05004125488104299500731A928380FF803DFBA0",
            INIT_RAM_2E => X"7C2EB9F5019B08800B002480260A1E1E068A8800010800010422090405908E94",
            INIT_RAM_2F => X"09018882CF4DDD0AA00021921BC4F5F86CBD8640F02489367FC00E00D2035000",
            INIT_RAM_30 => X"72C4771BC9E49462862410E05D123DA12AE1210980D006098394182763238224",
            INIT_RAM_31 => X"12484E950CC56BC2074E6383E8B04042283360C798A6D05587A80E3008028803",
            INIT_RAM_32 => X"EEBBEE57FADD8755954D598EEB4DD9A229110490C11A160050C0C240927D145F",
            INIT_RAM_33 => X"D1F0BCB00BFA88434FB28002164BAA0B6AA38801D622A4EB12B96B77DDA97FBB",
            INIT_RAM_34 => X"70C0C0AE65C005A47A90C935280105DC3D20488A6E0F1AC910FBDB1BCC2AA598",
            INIT_RAM_35 => X"531891B58D18DC176E107DD04E53D9EECBD895A915AD410510A830F00CA0CB67",
            INIT_RAM_36 => X"331F88D861240142CC0460CC6ED6BFC44D54D440A0460CC6E96BFC44D54D440A",
            INIT_RAM_37 => X"02E2221C980ACE30B33E40480610B0D0E3177C648495041100558E19667242D2",
            INIT_RAM_38 => X"1F18C040C1001C8BB1B16C102500019504905060BCE070204B89602430ADB088",
            INIT_RAM_39 => X"151F4BD011085515625D20155151515155555154107060A80203913071B8B134",
            INIT_RAM_3A => X"011D67811B0620585948DC092048CE307904C8B38052CD9F350C017047BAAB50",
            INIT_RAM_3B => X"09F34322045180C00B394151073201301238A684BC948C8902DA026041D2B1AA",
            INIT_RAM_3C => X"1DE4501D9A0FE6CFFD1420848E9DA29E29BAE7F0CE6004C0AA82011FB7D30029",
            INIT_RAM_3D => X"39B8701301A7180496217FDF81BCB510C2C067684008231D408A3D8C61150410",
            INIT_RAM_3E => X"7114A424525184619D891CA1596018620788140586C43189489624DC2B22684B",
            INIT_RAM_3F => X"01FEBFA30BE75228A800DE41F91E02F8C2F6C9122C24FCFCFB6342A01037601C"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"80D0C632F4DC8D192D59F1440612A3B1C24DF7E684CE802D4C39552000030481",
            INIT_RAM_02 => X"28E34CCE5D9DE4890B6F301809E388D551CCFFB836694494DF4FCBF4DA6FA65E",
            INIT_RAM_03 => X"2791B19772426BBB924924554010484D33DD8884DAAAAAF6FF50A78DFD9335A5",
            INIT_RAM_04 => X"5A1290609EF0A40CE5977F5B7E49212C9BB6F7F9572712878A4290CA2DD3FFF3",
            INIT_RAM_05 => X"48354A52141484916CAC00551A1B598D0BA0E5310A22890AA2D02114C96458A6",
            INIT_RAM_06 => X"04924926789272E52E9A08F142019031CA132084320637284C001C0A39032181",
            INIT_RAM_07 => X"689B51F90940C180C4C0B31254924922060ACF030483CDEC9F22C848CFE12C98",
            INIT_RAM_08 => X"EADE3D24C3F6236D701F3F07211301B72F74360E318C2043126447B8D928DDA5",
            INIT_RAM_09 => X"E3E73058FD3C8D9752512CF5B49C2F780F3FF8C57C57E872F3F539C9A4D8C09A",
            INIT_RAM_0A => X"2E9B61507DD55D9E5D90924932FB483AF68BDEDFE1F4DADE18DF0CE766C3C419",
            INIT_RAM_0B => X"6671E0E8300BFE6FDF674D224391D63E4080DF6830DACD930E713322333C6FBE",
            INIT_RAM_0C => X"4A0E4DAE263613E7D50A461A8C2EE4024267A1C4B4068B44D9211D54C25909A6",
            INIT_RAM_0D => X"1E60616364F44D3ECC1B46938D267BC302626135DC9A67B1611B883C0D319707",
            INIT_RAM_0E => X"2B10E73059C78DFFAE3ECC6F92699A7677672238DE498CE66178C7C5B3156333",
            INIT_RAM_0F => X"F3320809880A84C7C9C460C4CB805514450BD5DB59C595E514090A0184C69B04",
            INIT_RAM_10 => X"D8C201A0C15297E97D6410005BEF717A74A4F3FE3EE1440D414085500045B2B3",
            INIT_RAM_11 => X"F06545410236630034D2402106518098203DF7057481D60C07514E2106DD23DE",
            INIT_RAM_12 => X"48F29D50182002800AD22C3508E044434826434519412102C4992682980039D5",
            INIT_RAM_13 => X"D053A442B0C402804440A1E34682B840843027E42610E4023612B3153B188B10",
            INIT_RAM_14 => X"3502AEAA6C0108888224A962935D715B15502968AA82A2A56C4C20F4ECCA101E",
            INIT_RAM_15 => X"D45EA51C33CDF266261ACAC762E6B133861052380CF092F74B1602AB46EA32AA",
            INIT_RAM_16 => X"1440177620303B03302C674BAC89FB86AAA20904D4848C976A94A3AA21739518",
            INIT_RAM_17 => X"5294C1144AD6C9240234DA3AC9A325B707FC10671859246A83E513B2AED4711B",
            INIT_RAM_18 => X"29A1243408A0E9E68405045448190F80AA551650095493EE999C460E12066811",
            INIT_RAM_19 => X"F0B1AFC042898CF0CAAAA2322B96923E69307269A504AE098E164D8351255550",
            INIT_RAM_1A => X"DF1231DCB3030A520518AA01408A8A2006820286DE922128020020B438B006F0",
            INIT_RAM_1B => X"8A0843E9EA253C6BA7259280556B71785100E3E05ED87D5900941C12636B6383",
            INIT_RAM_1C => X"0088A342BD9140BC6D6D6B1CB1702A0AA9821A1DC946AF635360056D447D10A2",
            INIT_RAM_1D => X"344AA2C887707B6406AE229A271303C51120176063663108C7C2201F07FFC002",
            INIT_RAM_1E => X"A1CE610800970848FFDB891242A1623526662E01516D249984CF6D24ED64F693",
            INIT_RAM_1F => X"207100001B8E550E15560F1C35D0AA84370438C484147073F3FAE4F6D8879E30",
            INIT_RAM_20 => X"0129C093ADB6B182A00230AAA066739E346EA504545080CC82C040431143201B",
            INIT_RAM_21 => X"AEBBC35EB2320A8460644900898AED2031455464E8C48499E48932402D0E6880",
            INIT_RAM_22 => X"72823500044CEA3F0929421084C20551655A925944F4D42B4542225340864554",
            INIT_RAM_23 => X"2AD5542A1401F0CBBBBA5BC16C92B5B62C95916E9B0F5862E6D263B41C01212A",
            INIT_RAM_24 => X"9490A1771448824044555200A1AA82022226054142F0708044462050C952AD12",
            INIT_RAM_25 => X"C00E976BBB8A85014010316E923A188808628D085158AAA882A82ED4A4080A29",
            INIT_RAM_26 => X"140CE2482294E5BE7D01D1E963067A98C578A5F8C9F14E80910A857507BB88A0",
            INIT_RAM_27 => X"8A14E081CA0B40A9286A323940020000412602400499E11541C0604A2D557110",
            INIT_RAM_28 => X"05CB00008088822AE30CBAE310515394A09F14441102478822AB3106081031C0",
            INIT_RAM_29 => X"8A96B450E00000208D7CB294212007525CA9D6264AB9F30900000E2336036000",
            INIT_RAM_2A => X"15C0220977F36411145202AA06C82A086AD5613E89801281997E60A927161146",
            INIT_RAM_2B => X"F0EBE105E091A4200C007281F534272B90A95222B012AD66B182A0019564B529",
            INIT_RAM_2C => X"3BD26E3453363E8B4158A9158AB5A841DDD806E06075A10AF1342830952443B0",
            INIT_RAM_2D => X"3F8FFCC46F5E387813A5F834DE77882A5689652E74C0D270E1CF24A086FBFECE",
            INIT_RAM_2E => X"17BB3518F0C2BD8E7290E562A0699F1F0E0A4E0095C533DF4A7D6AE73745E4F9",
            INIT_RAM_2F => X"9A3887969A18857A4E3B0E406AA3AD51C5AB8CCCA4CC98A094163A63A186D604",
            INIT_RAM_30 => X"7CE6B15DCA3454811E3923A13287510ED701738E98070C28338C28619028054C",
            INIT_RAM_31 => X"0A602B5E88840C2D088084410210706004836E98420EA380C001E291B9BB101E",
            INIT_RAM_32 => X"554455E005229B8822000100404881030198A3EB9EAD72B5CAAA9140512884D4",
            INIT_RAM_33 => X"A224909649E085232E3046E173493580550111008901A644B455CEAA22380044",
            INIT_RAM_34 => X"991129C70321500822487418982B3170E04212000828C726810C24E43180BA2A",
            INIT_RAM_35 => X"00CBCE4070E526B05E22002208810201108E40F0C2101BE0CE03040450760691",
            INIT_RAM_36 => X"6A812457D0A7F50008A88E140140400280BE3F3F4A88E100100400280BE3F3F4",
            INIT_RAM_37 => X"B4101D518206333B634BCC5C66C1209041A51482922ABAE211AA4124D5CA080A",
            INIT_RAM_38 => X"7435AE01B1AC0D3390D2D686BB26ED29F9260F3603338B8E1208594D280824F3",
            INIT_RAM_39 => X"206E5F2E447E7777157A30204042C0C06040404129AAE4FD9C2EC471F5A82D77",
            INIT_RAM_3A => X"6BADEF984704EA310032F9092458853A7E4DE9A6E86DD0B08AC302028CC4548D",
            INIT_RAM_3B => X"200813B322AECF2E099477727FF211301B148BF6A2742309924CB4384DD191A8",
            INIT_RAM_3C => X"3CC1A90DDBC6828AA800E7315A0C801E5D900004D41DC0CABAE394608008BBBB",
            INIT_RAM_3D => X"EE6B29BE7FBD9756D660D537C9AAF59CE992636CE2BB3F1243D27B0DA3E72663",
            INIT_RAM_3E => X"372434234048AE2ABD096C02704D52225A29EA4B14DE379D488421080C004598",
            INIT_RAM_3F => X"642EC934401DD01BFF9BD404A0B5F29AF42487BA68DB0103776726C332732008"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"328004990002F148940488B22CA1952124824208488008728200000201E01002",
            INIT_RAM_02 => X"0690810106C5A2C0424A20525010420088198404A8D1A9D08121B2016CB48800",
            INIT_RAM_03 => X"0B0004200010100004020CD542380202448908A124104024812F04290505C3F8",
            INIT_RAM_04 => X"284688323DFBF64004121000219129010C4090008102A0285414051089228217",
            INIT_RAM_05 => X"03B0425A1024D240AC240006026840069C23B435432AA94288152A5125154AA1",
            INIT_RAM_06 => X"8B124A5878269018C020828884EB9040240013097208009000000550A6D7CB82",
            INIT_RAM_07 => X"03E4C5FDFCF8087808173620D00C492188112472E57B12E55A3CDACF1A166520",
            INIT_RAM_08 => X"9110241282040A4A491124924984D8C4B15E242A250840B02222212400148012",
            INIT_RAM_09 => X"1A122110A492400405044800000351800CD59660520506472A2E5D209280BB94",
            INIT_RAM_0A => X"09A25EBC496001300005200040821CCC09001490931294921689048424222196",
            INIT_RAM_0B => X"0341008220C00000014E885A928534A4604892401290490A63164811DA214304",
            INIT_RAM_0C => X"A56929114948A04508A861D04912430104209021CA895CAD6018D0000610500C",
            INIT_RAM_0D => X"0218920489420484062489250410500A00448AA550034524425014A408451415",
            INIT_RAM_0E => X"F1A0842915204920082420912440D081485C08A1249106914C0404B926404A12",
            INIT_RAM_0F => X"8C630324007B003268C9A1304CDC727025CA94DA6D8D350D6009EDF500130C28",
            INIT_RAM_10 => X"201EC20713209CCEC9251004F4006D01BAF5A2BA6BEBFABAFEBAEAEBBBEEBFFA",
            INIT_RAM_11 => X"0B90988C90C89885092CBAC2D1A48D609B88203B821A083060C3A055A9609821",
            INIT_RAM_12 => X"800A829601D5842C0700D15A6008198CA76B8CAC0228445C0A26607D255E43E1",
            INIT_RAM_13 => X"686D08B1B71ABF7B3566B3295423524484288420802C12014842408A0087243C",
            INIT_RAM_14 => X"3413CC004AB462222B18B3E68454401D1458E342099A4AA964AD5332ED1822C3",
            INIT_RAM_15 => X"659B383646ED81991047E4490228E66670C68D0684A08CE688248EB162BC6807",
            INIT_RAM_16 => X"082CD9B672A686244D6888AA28A858540008A4D0000946F99749F8FA0153F7E9",
            INIT_RAM_17 => X"5B5BE794AAD4018448914A8A89209097304192337998F8A8A1572D8EB37832DA",
            INIT_RAM_18 => X"AAA2D1B4A208ED24D14155559AF668AAA55748D62051033A25533174585615D3",
            INIT_RAM_19 => X"84462995C6822C0E11C000126B924B09A4D85A28BC09ADA9364924B1A4514140",
            INIT_RAM_1A => X"C40BB37398AB14A5101200498105044F2010805B864A413298AAAA92EA0E8122",
            INIT_RAM_1B => X"0A0850AA69822069A511000055689325533C494908498DE003D9218488D5E672",
            INIT_RAM_1C => X"2251840EB53998A66735BC648DB6A80AB22A4186C8128848211B956DA428DAA2",
            INIT_RAM_1D => X"FBF2A62F6323C949B34C8401994130053632D7658A9A739C73A0200D0000A302",
            INIT_RAM_1E => X"449088C06098B49C00DA324006EC40948998A0A84000004111492402651C90CE",
            INIT_RAM_1F => X"144522435186486033AD11148D000A81188023800C8C45399B020026D9106C1A",
            INIT_RAM_20 => X"54680031B6DB18C015A89A0A004C6C0C9929C38894046C9288021B3A4D68A534",
            INIT_RAM_21 => X"3301306007070041860E016EB43B2EF11989415263108411800011299689A488",
            INIT_RAM_22 => X"2AA081018D8850480A31C05220108081403064E2E00019B8646CBC8013317640",
            INIT_RAM_23 => X"4554002A401908844444491404025290311A0804C0081220324025A48C061298",
            INIT_RAM_24 => X"1B6AD5999411282B48940186A2A008AD0381508E18C90A00CCDA6802A2040D4C",
            INIT_RAM_25 => X"89ABF8A8444C0000096968048005465AA22A60B0535202AB9ECDB33BDF8E6A68",
            INIT_RAM_26 => X"04483144209850010C99690964442680CD400425A81840844CCA4848D8CCC2A0",
            INIT_RAM_27 => X"B02181A082DA821234202020618050060091892502E965140809081A2D050523",
            INIT_RAM_28 => X"B8144555130991108208AAA200533137A001144000421000229B132648912544",
            INIT_RAM_29 => X"0318C653400000000E090A52108000041222440812085251E06B4AF1AE028AAA",
            INIT_RAM_2A => X"940022300008241000054011E90106382E1516020200300CE080C0131BB71180",
            INIT_RAM_2B => X"885848891172E1645100008051100C1863386710DA00E74398C2902485A0D631",
            INIT_RAM_2C => X"2A2E12100801529889C9E4F59A146D4A2226B134888EC00A0100049015002680",
            INIT_RAM_2D => X"3800096EA3460818034983544489843932541E8291282680C80C86AA5418FC57",
            INIT_RAM_2E => X"1DAB0FFE5086408028A8020049A01E1E1E0ECA0011A4236208451609C62080C3",
            INIT_RAM_2F => X"0880A00082088408120C12C848090403028112500202040B3E8390048498440F",
            INIT_RAM_30 => X"9DD76B397B7D89084280489205241182C50142200481100501524A9548102800",
            INIT_RAM_31 => X"CA172C509280282A4011C004554FCFDC505246042D76022030046AC2D4613022",
            INIT_RAM_32 => X"555555A555AA8422C89AA515159225325132E88B30A14B09A412648650826880",
            INIT_RAM_33 => X"A221212112DB36B369A513336512C020C40933848B4D2045A10736AAAAD95555",
            INIT_RAM_34 => X"122607998E3E0A51A52F46D25C418952220485259B186E300808000000006ADB",
            INIT_RAM_35 => X"048CA000000007253E43AABB992D315584A962A4C14A81180800C109A3933C11",
            INIT_RAM_36 => X"3307C51048A09DA52869B12CD5CD628A02717081469B12CD5CD628A027170814",
            INIT_RAM_37 => X"73208168900410A04A00C049052CCCE200F248B688A8CB64B0884125345A22D9",
            INIT_RAM_38 => X"8005298621B402C79068140EA09929A80260A0830026003480118838C8524110",
            INIT_RAM_39 => X"0E8B400E664455551408D02A2220242232323230628B40CD26F0C8A3E74C08A5",
            INIT_RAM_3A => X"65994F0802031AAC000C79104285685A93094D2668A4802000331CF033328945",
            INIT_RAM_3B => X"84046502180098000022889354E4984D8C2131A68458059244901920BDD18DA8",
            INIT_RAM_3C => X"2848AD86D282009AA84631D87D280809110C3000F84CA293EDB64240C0044CC4",
            INIT_RAM_3D => X"213043420125308EDC325514092B361696CC4A4B666C22130E9222C8C23644C8",
            INIT_RAM_3E => X"09307670E82008032D8030A0954350A66F44AB659E86610DEDDE765C4E08D76E",
            INIT_RAM_3F => X"65F6B6EC9110F44AB464D439F6D4035BAAA491B348900000424A0B028B3019C2"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"B87E179D3C83E31247F8DEA3A6A515299492184BA66C6DE59337765F37D35978",
            INIT_RAM_02 => X"167C20221CB5E718192BAE0941EF8C8A364DA08615FF55689D920B2765B48CF5",
            INIT_RAM_03 => X"07018035501003378201167F689A0200222D338434C34C26FC91B42D81040129",
            INIT_RAM_04 => X"88D7E29B3DD4D501E1874252791122209C64D3F880221004080300C6A4D23E06",
            INIT_RAM_05 => X"C6FD4739CCD3994F5E74EE5531CF26DCC83FE6D33D659629AAD56130F338C9A4",
            INIT_RAM_06 => X"BA00001033B270188006106310C32114869346206422921A051000641D06A328",
            INIT_RAM_07 => X"1F8020000800080008CE269079B8000F00442D9180E95CC45F7898DE158C4D1A",
            INIT_RAM_08 => X"C15DA6CCFBF5216B6491B45B2B122106505BB4ADA56B02228E666532008296DA",
            INIT_RAM_09 => X"D34FB55AB6412005B4910C08000D21800000054248049079676C5392DC82E116",
            INIT_RAM_0A => X"8DBB48B06147458E1204304100518F89015E96920A089E9B96F8D2B5949230DA",
            INIT_RAM_0B => X"C02D0C832F50000001230C1332C19E353724DA4DCAD36962CE5C6D5B13AC7178",
            INIT_RAM_0C => X"1085AFEA662C3B3C43D6D24CED5156BC919ECD9996E6D9688E5FDDD9318C5525",
            INIT_RAM_0D => X"FB0E9D316116164403A96794B6095861D3327BBCDB2D75B0794AD617CB24E653",
            INIT_RAM_0E => X"F31CE7395DBF6D8128B1DE6C152008B0236E8C1CF05C807DEEF61605D62D81DA",
            INIT_RAM_0F => X"286303B425BA290359FA3C18D96C9366850BBEB6C9E616078449B975A4D39CA5",
            INIT_RAM_10 => X"01200000000066817DF6ABABBFAEC23E050E4945404EEBA6FFFFBFFEBEBA4D15",
            INIT_RAM_11 => X"F000404000000000000000080000800000082001000000000041000000401000",
            INIT_RAM_12 => X"10012000A00040028009000010012010100010104410802000000000100001C0",
            INIT_RAM_13 => X"9EC4545667B0060822C46ED62E9CA210042307E0090100A000A0044004400080",
            INIT_RAM_14 => X"41EE0DAF49480C4EBF33648157BB7D64C98A109BB04BECA6BAB6A6C99785B05F",
            INIT_RAM_15 => X"2F511A1C07ED3B99400DF5A10446A23278E5B0F117EDD8B6839F90028D24ABB1",
            INIT_RAM_16 => X"7E6A0A99543070B24593489BEF490F89AAFAF934F4F28D2A902104507F72A8C4",
            INIT_RAM_17 => X"6B5B69B4FF34926B60FEA071B6CAD9D8CBA8644CC567E6B113CA8058158A59E7",
            INIT_RAM_18 => X"29A5487919E7770D679FD7D60D1217AFA7FC4C39A1D1DE38211907C367F9DE79",
            INIT_RAM_19 => X"52267497B12B37FD33C1447F2C76DB301AC6765943ECF936436DB6CA9A335F5F",
            INIT_RAM_1A => X"28FD5B2B19EDC421782DA5BABDB0B2C16F4C6DE47B24A0C341505149413C1F8B",
            INIT_RAM_1B => X"0F06437D1405AE90CE4AD0ADD7B7D8C579ABFDF88F8302EBBE218CA35CFA307E",
            INIT_RAM_1C => X"A8008020D2BA05D09F359D93029EE94BD32DB7927F87C66C23465D138E3A23A7",
            INIT_RAM_1D => X"6281A3818D9EB4706790C8088362CA2D18FAB9B74D42318C53F7F58FB7EF6AC1",
            INIT_RAM_1E => X"77B3BA395A634289FF6C0408D190DC3E589DF8B1B56DB688DBE492DF0A6F0126",
            INIT_RAM_1F => X"8087B06E6EE5F15ABE61C3DA2BD5F0282BDEED71A2E1A210ED1F1BDB6E5CC57F",
            INIT_RAM_20 => X"2015300A400022168A4020F0F3A060FA0653083C60F8EB0C8E0054832FCE7196",
            INIT_RAM_21 => X"C03A8A8180405ABE3590BF59C7C552440BE41E64B1986311E4D2448475FC176C",
            INIT_RAM_22 => X"C407FFB570F70EF45194962176042C16BBAB080016D48A458BDA20FB4D0A2835",
            INIT_RAM_23 => X"476141C0A1EBFD711112DA164B2652DF610A8A4B64D40C0B8B648ADB1768EDFB",
            INIT_RAM_24 => X"2911428AA188D443AC61E3F4050F1AF2375F54411FC27052222317FD03D3B068",
            INIT_RAM_25 => X"7CB648C3DCD1EFFAB68CDB6B6DC0B1243C514976A82441404070956A5BFC1505",
            INIT_RAM_26 => X"EB7255B8F969093E77F56A1FB677A5F720BD5A141F63A9E88010E5864754570F",
            INIT_RAM_27 => X"4E9DA445AC36FCE1EF1AAFEFE8A55A58AC26B4987F473AF5F3AE5B4994D7C2AE",
            INIT_RAM_28 => X"0F7D31119C344CCEBAEB249AFFAA832E5F9869B7DF3869AECC446A244C993377",
            INIT_RAM_29 => X"A94A52843FFBEFBEF110DDEFFFFAA6E3FDFFBBF7FFF16C1B606B5E3422052AAA",
            INIT_RAM_2A => X"A1AECCC3B00393CF7DF9FF9B74ACB0C37DA37FF79DE2ED9D3F26DEE02489ECA3",
            INIT_RAM_2B => X"E7D647FD8B060396DB6B6A29CA25AFD656B7497E86DE10D846343AAB70824294",
            INIT_RAM_2C => X"4445C18D77DAFF452F1D9A2345CD11A32320E3864C4417A0C672EFCEA03F725E",
            INIT_RAM_2D => X"2EC0D828CE9DBF76B2693C40DE8A5FC6C71FA3F4FEAAC1D486D5FD0FEAEF5A1F",
            INIT_RAM_2E => X"3C717B56F6B51BD6951D79F587FFFE0F170E020A852101EF823B4DCDC7D58C98",
            INIT_RAM_2F => X"F7FFFF2F19927FFFF7575EB4BE82FFD8776B2FEFADCFFBE643A7A7F079C7FA03",
            INIT_RAM_30 => X"18DEED0A5BD5B0FF0DDFA068C0186AC4D28184332F67AF5E3E7D3FE92FC7FFCF",
            INIT_RAM_31 => X"FCF3F8F1CD641C1CBFCE0D2D56B8404A828A4B1129550D007807BB05FE6F981E",
            INIT_RAM_32 => X"9999981DDBBB3A99367D9AF4D21D9AE7D39F3B9E61F3EFAB36D636FFE5AB7F34",
            INIT_RAM_33 => X"44C4989C49DC2A17D9E81556E309541FB9E68CB764A24F324DDE0199990DDDDD",
            INIT_RAM_34 => X"EBB7DB5AD7DB15ACCD51F9FEA5A28E481A7185DAE6F32FB4E8A7DB168955959C",
            INIT_RAM_35 => X"B329F5BA4E15DD6CFC80515574D6628BE71ED8E32A1053533B523CE99DACAEED",
            INIT_RAM_36 => X"2AB7DF2F8BCE0A02D71440CA0AA0DC119C787A0211440CE0AE0DC119C787A021",
            INIT_RAM_37 => X"9CAEDBA16217DA9461BD3A748516508A083BCFEF20C35591A233FBEF3A9CC3BD",
            INIT_RAM_38 => X"3CB5AF0CAB7544821466DEA7F2CC7B7E81E9A095E8B1C2679ECF5A6A6BAEEC74",
            INIT_RAM_39 => X"F4745FF099BA888863F0008C282A28282828282A31FE7D8A1DBBBB3BFF257B3F",
            INIT_RAM_3A => X"5F5FFBFC468628A44418BBDC48B18A7C5FA4DBEB5AEDB024443C5EFE73F25032",
            INIT_RAM_3B => X"DEFBC7D7A1A2C7090015919EDEE2912010A9E0ADD32333C95248D07AC1D07DAD",
            INIT_RAM_3C => X"207BAB46FDA231CFED1CE59B1D8808A81589ABE419FE286636D3C0AE6EBA044B",
            INIT_RAM_3D => X"E724694F83F71937BFE8F71EDB7C6C0E70ECFEF4F3443F8FBCFFE29BCBFC1AC4",
            INIT_RAM_3E => X"177BBD244AEC2B1E3FE47208BFC8F3B3CB59EAD3E7FD7FFBD4F73C0DCFA27506",
            INIT_RAM_3F => X"753248E9507D7CEEE485F49CB39E077E99BDF7D6FB120354E7F7B3135FBFFAC1"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0102651B802E24792832217C849153A14F6FA5FCC00298A048B00126004B3485",
            INIT_RAM_02 => X"2D0031935808003536CAA026A443A77CE1D9FA5C4DFFD9CF676A329A0007E20A",
            INIT_RAM_03 => X"93C1C63559090AAEC32192A89BC1212199795111AFBEBAF297016409297FE20E",
            INIT_RAM_04 => X"D0148B02B1B1A441A084494D8985C010CEDABFAC080048902108423092017CE1",
            INIT_RAM_05 => X"B22090942189F071498A1A8CE4F193260DE2FD40180C32C42AC549E1AE531202",
            INIT_RAM_06 => X"0B8006D910410B19C830293BC22D00523C487784A00A48F1210039224F5AE506",
            INIT_RAM_07 => X"6FFFDC0008780078003A0C6A5B6E0000BD314A89104E27586628318F02441820",
            INIT_RAM_08 => X"971229308A54044A58562B868B48A455AA40A40C2588E329BC8083A924188935",
            INIT_RAM_09 => X"0A32A910A9ACD2459644E8F90248807FF000066F52F46542DAC4794D228C9554",
            INIT_RAM_0A => X"082242C1553201840EC30000C904D9DC6541549172A6949410924884640AE017",
            INIT_RAM_0B => X"309142E8A14BFE6FDF35CC582281342E89C29F407091CD03EF6E90A592A85CEA",
            INIT_RAM_0C => X"C2124A3C78C6168A9C08CC20093EE646424BA14E80181C0B0103500444211A82",
            INIT_RAM_0D => X"2E9264CC58A1082F24981862088554C4800492281690552450219C4808122588",
            INIT_RAM_0E => X"68488425116DC95E8B2B998AE28C26CC8745C2430B8A210F41DCE5516338A422",
            INIT_RAM_0F => X"F550420858B6D02D40DB65546E1BEEA93E788793401A82483464DE0112564810",
            INIT_RAM_10 => X"FEDFFFFFFFFFF7FF7DBEBFBFAFBAFB2AEEBEBBFE7EBEAEBFFFFAFFFFEBFAFABF",
            INIT_RAM_11 => X"0FFFBFBFFFFFFFFFFFFFFFF7FFFF7FFFFFF7DFFEFFFFFFFFFFBEFFFFFFBFEFFF",
            INIT_RAM_12 => X"EFFEDFFF5FFFBFFD7FF6FFFFEFFEDFEFEFFFEFEF3BEF7FDFFFFFFFFFEFFFFE3F",
            INIT_RAM_13 => X"9A52269CD0BD43008610C29122B722448008A3C7C63EFF5FFF5FFBBFFBBFFF7F",
            INIT_RAM_14 => X"155B08AA4AA1084AA91FFD3371837564454143488B8AC30968E952F76DCA9A76",
            INIT_RAM_15 => X"89D77838752964EF1CDD6CAE008811C5F4D49FB209A48EA4811E0AAB437A5226",
            INIT_RAM_16 => X"080EE476C2A6BE057449AE938E48AAD6AAAAA484C4D6474011491B402A4A2245",
            INIT_RAM_17 => X"28C50614E0D249260E345A808DB5B5293189D8137898A8E221A8BF840824319A",
            INIT_RAM_18 => X"8202FCB4ABAE6DE6D658D5055A6D2BAAA7021E56ACD099D79CC0C5FC1A561C48",
            INIT_RAM_19 => X"B555EB40C4D28DFEF70000050484D9FF60AC5C41094410E93C136931775A1415",
            INIT_RAM_1A => X"C7D236A56EA24210200600C140C4C30986C204C5CE9341A8C9AAEB929A1A8F60",
            INIT_RAM_1B => X"000C402AEEA2226F3117A004854AF17D5309CB684079BD389BDC38D1B812E127",
            INIT_RAM_1C => X"227F1FDF6D31C0AEC14C722CB9E200083AA31A8FD344000A2050006D24288802",
            INIT_RAM_1D => X"9570541F07756D75664A09522601B142A5280361A05C00841242400317EF6383",
            INIT_RAM_1E => X"61F8401040DF285400D29F7A0447BA20BFFB6E00824924999DCE4926AF50F499",
            INIT_RAM_1F => X"A0730007192CD44216801F100A040022150020D40888706332CEA474D0C2FB1A",
            INIT_RAM_20 => X"2105108209248102A10220A0A30E0FD67E43628EE0506154000021525B40606D",
            INIT_RAM_21 => X"04B2A01C3030006D44FA1A4CA8A4915160EE1444C344008824C922433F2840C0",
            INIT_RAM_22 => X"50039C913A3300000084502142C201A30A20DA2A24600707031D70895B884EC1",
            INIT_RAM_23 => X"54C00040C00970D3333213D04E9021242489004E926E183564927536093583B0",
            INIT_RAM_24 => X"1641A35515DDC0038EF541C7A20A0AAE102D54698B77780000147B062A10105D",
            INIT_RAM_25 => X"DCB752AA230B20681B50404ED252209028410432596002805134EAB4A5C55B2D",
            INIT_RAM_26 => X"2616A1D06BA8A12E580388B34505F52E65AC0D4032E1C5A4CEFAE5AEEAAB84A0",
            INIT_RAM_27 => X"2222C101C015803B8DC1335AE306406C35B51B6D0613CDA011C23142B1007713",
            INIT_RAM_28 => X"007900000AD55554C30C30C32AAE83CA001A2082083035000030202040810385",
            INIT_RAM_29 => X"121084579FF9A69A603DF084210AA27746C8D1234480E519402100143E05EAAA",
            INIT_RAM_2A => X"154888A9C01D4208208A800034114514258237BE0AC0EE092DFE643A20092100",
            INIT_RAM_2B => X"80B2E0B356AD5259B62AD00060048412FA327034E00484421082B02021008421",
            INIT_RAM_2C => X"047084E093BF2C43E1B1DC2231A8082ABAB81D60A8A50200A0040C2480826310",
            INIT_RAM_2D => X"A90F5C444E1C38700289404086220D376C190320B40A7420A00B200A946B4289",
            INIT_RAM_2E => X"7DE1696A04C4398358302040E9EADE0F1E160208012000CC0402042BA428C0A2",
            INIT_RAM_2F => X"D8AD2A940000091A3621273A10220C0A810386C40C86AD028015A241318CD402",
            INIT_RAM_30 => X"72CFBDFE4B58BCCA1EAD03313FE53304C08152AF8603060C13D632B181092A04",
            INIT_RAM_31 => X"3B10EAD59EC420236ADE4505555F6F765052460C2F100800B0042AF72D1CA803",
            INIT_RAM_32 => X"555555655688C7AABBAEEDB5554EEDBAC0371ADB8BBB58496912CCD9DA823D60",
            INIT_RAM_33 => X"00836B61B6FA99C36FB544035DF6F4B5336EAC13326F31112445FA22AAF05511",
            INIT_RAM_34 => X"A931285C0C014E1D11205A124899226188813211124288A68A20400432D5C1F8",
            INIT_RAM_35 => X"B32F89AA320004E3FD03EB9AB588935CC239BAF32B5ACBCB77519C8DF18C3889",
            INIT_RAM_36 => X"F3369D6287B1428D6DC57F785C85AA888AC340BC1C57F785C85AA888AC340BC1",
            INIT_RAM_37 => X"F2302770C4174047444BC628C1C54059241E59A4CE0324102822DB6D601378D1",
            INIT_RAM_38 => X"80043325718C66B6C250100EC8A48D0278330004403081E40013396919110C19",
            INIT_RAM_39 => X"20A4402C221000101402300010119190101010131007E0ECB68CD3F334050DF3",
            INIT_RAM_3A => X"7BAC698A2A063A2F102EB19D42E52D53361B4927E8C9CA7ABBB003F03F907F2F",
            INIT_RAM_3B => X"3910E90A4B00C2072C47F7726578B48A45A57086A01801364DB45CD9BFFFBEAB",
            INIT_RAM_3C => X"16600DA79AD3E955137EF6F00E1E0018D5C44440F49D2131BCFB72019109DDD9",
            INIT_RAM_3D => X"FC6B28877F8B8774C62200070D032289059C6269C3551F021D926BC9A1E54C67",
            INIT_RAM_3E => X"9F21A458AC324F9F99AD680484020124D05D4369B4C6B18C47348DA088EF02B5",
            INIT_RAM_3F => X"F52E02525007081DAECBC03E04A00393F026C13249CAAAAB736B5F40B7747D66"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"8135427A4A642F7B1CC40B3D2EB95714EDB4CED9D55639AAC28AAB0EAAE8742C",
            INIT_RAM_02 => X"2517D5D75372D72C2DAF3424AD94AE0AAA1DC5C84F00F442BB40B32E9B6EC23C",
            INIT_RAM_03 => X"B27152866B5B53315168BAAAAAAB6B6AAA9DE211BD34D2406A14460994E81144",
            INIT_RAM_04 => X"56B5CA4BBDF1EC0E45953616718DE334786CD0526B264E102148522AD2C2BF01",
            INIT_RAM_05 => X"3B7239DE731CE1739D90B1A45E74C56F5FC7B88EFB534CCE576A8AADD2EB3555",
            INIT_RAM_06 => X"AF924DBF7BE36969483B311BD2A63547BCFF77A5C6A8FEF3FD55702C475CEE2D",
            INIT_RAM_07 => X"7FFFFC0008040404040ABED8FA5E492FD975EAD9B14FAFFD796AFBDFD9AD7D9A",
            INIT_RAM_08 => X"DF1E192251A2A42E714E1D948F58E573152912A494AD816AA9D5D61D6D1CD936",
            INIT_RAM_09 => X"2A741D1A49A6D6D6273784F126DC80000F3C066E72E3C57AB8A56A4D36687DDC",
            INIT_RAM_0A => X"452320F528D0822101D2A249AB355CFE09D71ED332E6D65E589618D2E2A9C80B",
            INIT_RAM_0B => X"D484AAE2B550000258498DA80B41BC3CAA8A4E2AB0CA84A16B47B1E393386712",
            INIT_RAM_0C => X"E7120C7D718A21693A5D6D212564CB5740E5B24EAAB54EAE832B4AACD6AB408C",
            INIT_RAM_0D => X"56BA76DAB54B5D5D6E9AB1C55DAA7DC42AAAA772BCD067346523184CA5520388",
            INIT_RAM_0E => X"7A42D6911BC284AD46142355D45520E088640A463751691200294291A7720473",
            INIT_RAM_0F => X"CF72B2A839B6813F459FF1DCEDBAEEFAAF5BCE9254AB8AEAAC3FDEABBB57EE91",
            INIT_RAM_10 => X"1124512422249B49A6DBEBBEEFAFFB3BBBFAFFBA6EABEFEAAAAABAFFABFFFBFA",
            INIT_RAM_11 => X"F89445449088844888A2410C0A44821041082089042041021041111088409111",
            INIT_RAM_12 => X"00100010008004000200101000100200002080004410892244924924909249E9",
            INIT_RAM_13 => X"EF5D4AA96A1FFFFBBBB75BFEF9738A74E72EE7E0000080008002000040008004",
            INIT_RAM_14 => X"4AB3ED556D777735553D7A9436EECA8FBABAC6477917EAF9E8D9BA62CD892AAA",
            INIT_RAM_15 => X"EFDF7CE9552DFEAB9C7F6EEFD7FF557515D0DD025E21DEC6CBBC7D58ACF6CDD5",
            INIT_RAM_16 => X"DDAABFF475744E2D7549AEAE79155D2C555555DA3A2DEE7FD7AD777F55FBB7ED",
            INIT_RAM_17 => X"D7BD6BAADF9DB7344EB6C5FE393648D5B26591F67091A8FFFEA7BD1FFFBD73D0",
            INIT_RAM_18 => X"D555D0B4D4516DA6CBAE2AFB1764745556FA5C5C3D2D55B625595D74522C5A5B",
            INIT_RAM_19 => X"87F76915E7DBA81EF7D5554B79DB254D12F9FB7DD8ADE55D344C96F32448AAAA",
            INIT_RAM_1A => X"8ED222A56EAA3FFF67BEFFDBBD7575EAEA3FEC8184277FA254411401D55D5362",
            INIT_RAM_1B => X"FFFDAAD648A6364D339592AC7ACFD932AB8A6C69E4C9B8FB9B993DD4B8B0E532",
            INIT_RAM_1C => X"2A00000027AB0767EEFBDEBEDBB2BFF7E2AA30949353D2AAABC017E82E480AFD",
            INIT_RAM_1D => X"FBFDF7459B23D0D9117CB782AE5B328FBCF20265AB3B394A52E66FCF2FFFAB3F",
            INIT_RAM_1E => X"E5B7FA2D5FD8629D499A3C7897579A9EBEFAC8A57DB6DB271561B6DC52BFDB8E",
            INIT_RAM_1F => X"8AE62D4B5BA4D946BFE8DFFEAEFCFFE6BB9F8D912EEDC5FFDA365BA699D4FD33",
            INIT_RAM_20 => X"DF782FB8FFFFBFF57FBE8F5F51EE6E32BF35FBEABEAAC1146B79E5575E6AC564",
            INIT_RAM_21 => X"BF8802FDF3F3DEED159EB85D627BE77DFAABEA896754E711DB46D48573BDF388",
            INIT_RAM_22 => X"EFD56AD15FCC9AED5D7BAFDEE5CE6FBCF72BCCFAFBBEBD7EEEBFFEFAB9B7B6BF",
            INIT_RAM_23 => X"57FFEABF9FEB918EEEECED95B46FFEDCEBFFFBB4CDC9F9B7B36DB7A67D24DF72",
            INIT_RAM_24 => X"2ECE7CCEAB157F7F8AAABBC555F5D55CFA52AAAAD440F5FAEEF3577EABF7EE5D",
            INIT_RAM_25 => X"8543ACD5FEDD27E9FB4D9BB48DEFFFFBD73EF8FCAA8FFD7DD7555DAC63CF7550",
            INIT_RAM_26 => X"E45A55CAE98D5ED1ADFF7A7B655F2DA6AA14FCBDFA1ACB8AAAA52A0AA976545F",
            INIT_RAM_27 => X"CA1EF5F4BF5DFFE39DBEEF6D74BC53C2E44AB092FEFF691FEA894ADD46FFC72F",
            INIT_RAM_28 => X"8F787555D62DDDDFBEFBEFBED553B97AAA8DDF7DF7CF74FFFFDD73A74E9D3D37",
            INIT_RAM_29 => X"EDEF7AAB600659659399DBDEF7B556676E6D9BB66EDF3E1D11A525495009C002",
            INIT_RAM_2A => X"AB377767981BBFFFFFFAEA922D3DF7DF7F9E63A6DD817EDC39A05BE3C031DEFB",
            INIT_RAM_2B => X"E59F4EEEDDBB797A7D554FFD5FBE2EDF7BBDFF63FEFB7B1DEF7567AEDEFB7BDE",
            INIT_RAM_2C => X"486257DF791324C987F1F83EEAD9254ABABA9554AEADD5FF8FEBFCFB9D5DE3FB",
            INIT_RAM_2D => X"B3FF09C4F9F3E7C7BBADDC7E9CA0DDBE7C1DA3B7E6AEC77EE55933F59A18D76A",
            INIT_RAM_2E => X"F004E2002BB7491E31B9E1C78EED9E1F1F9FC21295A5326CCA5E476BB7EEBEEB",
            INIT_RAM_2F => X"93D9B63CFFDFFDF3FE73905EFBE8F9FBFF3E3C9CF46CFDBEFFA5C647E7139E10",
            INIT_RAM_30 => X"C520C0D41DCF186D74F9AEF0FFFCAF2BC8C0CE623C773E7CB26E1B732787B76C",
            INIT_RAM_31 => X"BB3AEDDB848175766555EAAAACBACACAAAAB6ED3FFF55F7562AEF72B2D5BB85D",
            INIT_RAM_32 => X"EEEEFFB6ECFFDC55D575590AAB1559356ABA4FBA6FA74F793D726FCDDBD77D8A",
            INIT_RAM_33 => X"55D6DE4564D22F776D32D7F74B2DCBABEEABBBA5DE2B32EF23BFB7FF77D13BFF",
            INIT_RAM_34 => X"0266421C8E464B4D05303A0A6DDF44899DD2648406175FF62B610009067EC5F1",
            INIT_RAM_35 => X"F67D1D3E07004C1FFDFEBEDBD5A03BF6877FAFA77DEFD11FB1FAC9D985893C23",
            INIT_RAM_36 => X"FC1FDD1D6FB2AAAAC8D571FCF6CF3FFDDFF9F9C2AD571FCF6CF3FFDDFF9F9C2A",
            INIT_RAM_37 => X"F772AF65CA02644924588841455550C3655248E6CE967195AB77CF3D27FB7A99",
            INIT_RAM_38 => X"C0AD7DAF63962FB7D6E5BEECB4E95994026040409044202C5555A83958405950",
            INIT_RAM_39 => X"911A0F108028B3A277FDC33282828082828282814953EDDDBCDDD5F3F74559F5",
            INIT_RAM_3A => X"4B9DEBBD5702FABF557EFB146AF5AE733F36ED366C9286E5C3C0140EE62AC4C1",
            INIT_RAM_3B => X"E5557B9F2E4110812547FFF35C68F58E5739B9AC8AAAAB2D5B6ABCBB7FFFFEA9",
            INIT_RAM_3C => X"3AC759AE9B974A555556B46AAC32AABDD95D75541928A9376DBE66D5D559F77B",
            INIT_RAM_3D => X"E2B603C301B1299ECEF22A8ED995F79D179EE76DC7773F172F9A62D9C8F454EF",
            INIT_RAM_3E => X"A932F656AABAAAAB092472AC8EAAAA75556D16631EDE77BCE55E55552D2AAFBD",
            INIT_RAM_3F => X"E5390F7FD17FF2AEE76DCABD55A0063BF5768F3B4CB45454EF6F6DD2EBF7FD6E"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM_apple2
