--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.10.03 (64-bit)
--Part Number: GW5AT-LV60PG484AC1/I0
--Device: GW5AT-60
--Device Version: B
--Created Time: Thu Jun 12 13:38:05 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_SDPB_8k is
    port (
        dout: out std_logic_vector(7 downto 0);
        clka: in std_logic;
        cea: in std_logic;
        clkb: in std_logic;
        ceb: in std_logic;
        oce: in std_logic;
        reset: in std_logic;
        ada: in std_logic_vector(12 downto 0);
        din: in std_logic_vector(7 downto 0);
        adb: in std_logic_vector(12 downto 0)
    );
end Gowin_SDPB_8k;

architecture Behavioral of Gowin_SDPB_8k is

    signal sdpb_inst_0_dout_w: std_logic_vector(29 downto 0);
    signal sdpb_inst_1_dout_w: std_logic_vector(29 downto 0);
    signal sdpb_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal sdpb_inst_3_dout_w: std_logic_vector(29 downto 0);
    signal gw_gnd: std_logic;
    signal sdpb_inst_0_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_0_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_0_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_0_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_0_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_1_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_1_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_1_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_1_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_1_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_2_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_2_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_2_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_2_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_2_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_3_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_3_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_3_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_3_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_3_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_3_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component SDPB
        generic (
            READ_MODE: in bit := '0';
            BIT_WIDTH_0: in integer :=16;
            BIT_WIDTH_1: in integer :=16;
            BLK_SEL_0: in bit_vector := "000";
            BLK_SEL_1: in bit_vector := "000";
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLKA: in std_logic;
            CEA: in std_logic;
            CLKB: in std_logic;
            CEB: in std_logic;
            OCE: in std_logic;
            RESET: in std_logic;
            BLKSELA: in std_logic_vector(2 downto 0);
            BLKSELB: in std_logic_vector(2 downto 0);
            ADA: in std_logic_vector(13 downto 0);
            DI: in std_logic_vector(31 downto 0);
            ADB: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    sdpb_inst_0_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_0_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_0_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_0_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(1 downto 0);
    sdpb_inst_0_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(1 downto 0) <= sdpb_inst_0_DO_o(1 downto 0) ;
    sdpb_inst_0_dout_w(29 downto 0) <= sdpb_inst_0_DO_o(31 downto 2) ;
    sdpb_inst_1_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_1_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_1_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_1_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(3 downto 2);
    sdpb_inst_1_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(3 downto 2) <= sdpb_inst_1_DO_o(1 downto 0) ;
    sdpb_inst_1_dout_w(29 downto 0) <= sdpb_inst_1_DO_o(31 downto 2) ;
    sdpb_inst_2_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_2_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_2_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_2_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(5 downto 4);
    sdpb_inst_2_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(5 downto 4) <= sdpb_inst_2_DO_o(1 downto 0) ;
    sdpb_inst_2_dout_w(29 downto 0) <= sdpb_inst_2_DO_o(31 downto 2) ;
    sdpb_inst_3_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_3_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_3_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_3_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(7 downto 6);
    sdpb_inst_3_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(7 downto 6) <= sdpb_inst_3_DO_o(1 downto 0) ;
    sdpb_inst_3_dout_w(29 downto 0) <= sdpb_inst_3_DO_o(31 downto 2) ;

    sdpb_inst_0: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"0AA82AAA2AAA2AAA2AAA080000002AAA0AA82AAA2AAA2AAA0AA82AAA2AA00AA8",
            INIT_RAM_01 => X"C0000200200200082AAA2802000A280A2AAA02AA0AAA000208282AAA0AA82AAA",
            INIT_RAM_02 => X"080000000080000000800808000002A000000A28080A08202080000000000000",
            INIT_RAM_03 => X"00080000022000800000000020280A2800020AA0082A02800802280800000AA8",
            INIT_RAM_04 => X"3F7C0000D1FFFFFCFF9FF6FF7FFFFD1FFCCF4E9F02C0FDBF1FF4555F5A9F501F",
            INIT_RAM_05 => X"AAAA3FFCFCCF3FFCFD1FFFFFCFCFCAA766669999FF3F2AAAFF3FFC7FFD3F3F3F",
            INIT_RAM_06 => X"0A802AA02AA000002AAA200000002AAA028000800A800A800A802AAA08000000",
            INIT_RAM_07 => X"08880008200200000080202002A020202AA002A00AA0002020802AA00280AAA0",
            INIT_RAM_08 => X"F557D555D555D555D555F7FFFFFFD555F557D555D555D555F557D555D55FF557",
            INIT_RAM_09 => X"3FFFFDFFDFFDFFF7D555D7FDFFF5D7F5D555FD55F555FFFDF7D7D555F557D555",
            INIT_RAM_0A => X"F7FFFFFFFF7FFFFFFF7FF7F7FFFFFD5FFFFFF5D7F7F5F7DFDF7FFFFFFFFFFFFF",
            INIT_RAM_0B => X"FFF7FFFFFDDFFF7FFFFFFFFFDFD7F5D7FFFDF55FF7D5FD7FF7FDD7F7FFFFF557",
            INIT_RAM_0C => X"F557D555D555D555D555F7FFFFFFD555F557D555D555D555F557D555D55FF557",
            INIT_RAM_0D => X"3FFFFDFFDFFDFFF7D555D7FDFFF5D7F5D555FD55F555FFFDF7D7D555F557D555",
            INIT_RAM_0E => X"F57FD55FD55FFFFFD555DFFFFFFFD555FD7FFF7FF57FF57FF57FD555F7FFFFFF",
            INIT_RAM_0F => X"F777FFF7DFFDFFFFFF7FDFDFFD5FDFDFD55FFD5FF55FFFDFDF7FD55FFD7F555F",
            INIT_RAM_10 => X"F000F515FA2AFF3FF040F555FA6AFF7FF080F595FAAAFFBFF0C0F5D5FAEAFFFF",
            INIT_RAM_11 => X"E000E515EA2AEF3FE040E555EA6AEF7FE080E595EAAAEFBFE0C0E5D5EAEAEFFF",
            INIT_RAM_12 => X"D000D515DA2ADF3FD040D555DA6ADF7FD080D595DAAADFBFD0C0D5D5DAEADFFF",
            INIT_RAM_13 => X"C000C515CA2ACF3FC040C555CA6ACF7FC080C595CAAACFBFC0C0C5D5CAEACFFF",
            INIT_RAM_14 => X"B000B515BA2ABF3FB040B555BA6ABF7FB080B595BAAABFBFB0C0B5D5BAEABFFF",
            INIT_RAM_15 => X"A000A515AA2AAF3FA040A555AA6AAF7FA080A595AAAAAFBFA0C0A5D5AAEAAFFF",
            INIT_RAM_16 => X"900095159A2A9F3F904095559A6A9F7F908095959AAA9FBF90C095D59AEA9FFF",
            INIT_RAM_17 => X"800085158A2A8F3F804085558A6A8F7F808085958AAA8FBF80C085D58AEA8FFF",
            INIT_RAM_18 => X"700075157A2A7F3F704075557A6A7F7F708075957AAA7FBF70C075D57AEA7FFF",
            INIT_RAM_19 => X"600065156A2A6F3F604065556A6A6F7F608065956AAA6FBF60C065D56AEA6FFF",
            INIT_RAM_1A => X"500055155A2A5F3F504055555A6A5F7F508055955AAA5FBF50C055D55AEA5FFF",
            INIT_RAM_1B => X"400045154A2A4F3F404045554A6A4F7F408045954AAA4FBF40C045D54AEA4FFF",
            INIT_RAM_1C => X"300035153A2A3F3F304035553A6A3F7F308035953AAA3FBF30C035D53AEA3FFF",
            INIT_RAM_1D => X"200025152A2A2F3F204025552A6A2F7F208025952AAA2FBF20C025D52AEA2FFF",
            INIT_RAM_1E => X"100015151A2A1F3F104015551A6A1F7F108015951AAA1FBF10C015D51AEA1FFF",
            INIT_RAM_1F => X"000005150A2A0F3F004005550A6A0F7F008005950AAA0FBF00C005D50AEA0FFF",
            INIT_RAM_20 => X"0AA82AAA2AAA2AAA2AAA080000002AAA0AA82AAA2AAA2AAA0AA82AAA2AA00AA8",
            INIT_RAM_21 => X"C0000200200200082AAA2802000A280A2AAA02AA0AAA000208282AAA0AA82AAA",
            INIT_RAM_22 => X"080000000080000000800808000002A000000A28080A08200220000000000000",
            INIT_RAM_23 => X"00080000022000800000000020280A2800020AA0082A02800802280800000AA8",
            INIT_RAM_24 => X"3F7C0000D1FFFFFCFF9FF6FF7FFFFD1FFCCF4E9F02C0FDBF1FF4555F5A9F501F",
            INIT_RAM_25 => X"AAAA3FFCFCCF3FFCFD1FFFFFCFCFCAA766669999FF3F2AAAFF3FFC7FFD3F3F3F",
            INIT_RAM_26 => X"0A802AA02AA000002AAA200000002AAA028000800A800A800A802AAA08000000",
            INIT_RAM_27 => X"08880008200200000080202002A020202AA002A00AA0002020802AA00280AAA0",
            INIT_RAM_28 => X"F557D555D555D555D555F7FFFFFFD555F557D555D555D555F557D555D55FF557",
            INIT_RAM_29 => X"3FFFFDFFDFFDFFF7D555D7FDFFF5D7F5D555FD55F555FFFDF7D7D555F557D555",
            INIT_RAM_2A => X"F7FFFFFFFF7FFFFFFF7FF7F7FFFFFD5FFFFFF5D7F7F5F7DFFDDFFFFFFFFFFFFF",
            INIT_RAM_2B => X"FFF7FFFFFDDFFF7FFFFFFFFFDFD7F5D7FFFDF55FF7D5FD7FF7FDD7F7FFFFF557",
            INIT_RAM_2C => X"F557D555D555D555D555F7FFFFFFD555F557D555D555D555F557D555D55FF557",
            INIT_RAM_2D => X"3FFFFDFFDFFDFFF7D555D7FDFFF5D7F5D555FD55F555FFFDF7D7D555F557D555",
            INIT_RAM_2E => X"F57FD55FD55FFFFFD555DFFFFFFFD555FD7FFF7FF57FF57FF57FD555F7FFFFFF",
            INIT_RAM_2F => X"F777FFF7DFFDFFFFFF7FDFDFFD5FDFDFD55FFD5FF55FFFDFDF7FD55FFD7F555F",
            INIT_RAM_30 => X"F000F515FA2AFF3FF040F555FA6AFF7FF080F595FAAAFFBFF0C0F5D5FAEAFFFF",
            INIT_RAM_31 => X"E000E515EA2AEF3FE040E555EA6AEF7FE080E595EAAAEFBFE0C0E5D5EAEAEFFF",
            INIT_RAM_32 => X"D000D515DA2ADF3FD040D555DA6ADF7FD080D595DAAADFBFD0C0D5D5DAEADFFF",
            INIT_RAM_33 => X"C000C515CA2ACF3FC040C555CA6ACF7FC080C595CAAACFBFC0C0C5D5CAEACFFF",
            INIT_RAM_34 => X"B000B515BA2ABF3FB040B555BA6ABF7FB080B595BAAABFBFB0C0B5D5BAEABFFF",
            INIT_RAM_35 => X"A000A515AA2AAF3FA040A555AA6AAF7FA080A595AAAAAFBFA0C0A5D5AAEAAFFF",
            INIT_RAM_36 => X"900095159A2A9F3F904095559A6A9F7F908095959AAA9FBF90C095D59AEA9FFF",
            INIT_RAM_37 => X"800085158A2A8F3F804085558A6A8F7F808085958AAA8FBF80C085D58AEA8FFF",
            INIT_RAM_38 => X"700075157A2A7F3F704075557A6A7F7F708075957AAA7FBF70C075D57AEA7FFF",
            INIT_RAM_39 => X"600065156A2A6F3F604065556A6A6F7F608065956AAA6FBF60C065D56AEA6FFF",
            INIT_RAM_3A => X"500055155A2A5F3F504055555A6A5F7F508055955AAA5FBF50C055D55AEA5FFF",
            INIT_RAM_3B => X"400045154A2A4F3F404045554A6A4F7F408045954AAA4FBF40C045D54AEA4FFF",
            INIT_RAM_3C => X"300035153A2A3F3F304035553A6A3F7F308035953AAA3FBF30C035D53AEA3FFF",
            INIT_RAM_3D => X"200025152A2A2F3F204025552A6A2F7F208025952AAA2FBF20C025D52AEA2FFF",
            INIT_RAM_3E => X"100015151A2A1F3F104015551A6A1F7F108015951AAA1FBF10C015D51AEA1FFF",
            INIT_RAM_3F => X"000005150A2A0F3F004005550A6A0F7F008005950AAA0FBF00C005D50AEA0FFF"
        )
        port map (
            DO => sdpb_inst_0_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_0_BLKSELA_i,
            BLKSELB => sdpb_inst_0_BLKSELB_i,
            ADA => sdpb_inst_0_ADA_i,
            DI => sdpb_inst_0_DI_i,
            ADB => sdpb_inst_0_ADB_i
        );

    sdpb_inst_1: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"3003009000A43000026030003AAB00C0300300C330C33003300330C3030632A3",
            INIT_RAM_01 => X"C000006030030090355731832A9001900680240030002AAB30C302C3320300C3",
            INIT_RAM_02 => X"0180200000C01A000AE82BBA20022406002A326901852EEE25D6001522AA0000",
            INIT_RAM_03 => X"22831809033009181A20022030C330C3158330C630330318308331833AAE3183",
            INIT_RAM_04 => X"34070000A2BFFFFC555145557FFFDB39D2E7CDCF1600E9FF196CE0BF9FE78027",
            INIT_RAM_05 => X"FFFF3C3CEAEA3FFCD001FFFFCFCFCFF366669999DF3D3FFFFF3FD407D0176002",
            INIT_RAM_06 => X"303000300A903AAB0300C0203AB20030CC3015D6333030303030303033300009",
            INIT_RAM_07 => X"0998000B3A2BAAAA2F7E3630CC0006401A00240030002575333000600C300C30",
            INIT_RAM_08 => X"CFFCFF6FFF5BCFFFFD9FCFFFC554FF3FCFFCFF3CCF3CCFFCCFFCCF3CFCF9CD5C",
            INIT_RAM_09 => X"3FFFFF9FCFFCFF6FCAA8CE7CD56FFE6FF97FDBFFCFFFD554CF3CFD3CCDFCFF3C",
            INIT_RAM_0A => X"FE7FDFFFFF3FE5FFF517D445DFFDDBF9FFD5CD96FE7AD111DA29FFEADD55FFFF",
            INIT_RAM_0B => X"DD7CE7F6FCCFF6E7E5DFFDDFCF3CCF3CEA7CCF39CFCCFCE7CF7CCE7CC551CE7C",
            INIT_RAM_0C => X"CFFCFF6FFF5BCFFFFD9FCFFFC554FF3FCFFCFF3CCF3CCFFCCFFCCF3CFCF9CD5C",
            INIT_RAM_0D => X"3FFFFF9FCFFCFF6FCAA8CE7CD56FFE6FF97FDBFFCFFFD554CF3CFD3CCDFCFF3C",
            INIT_RAM_0E => X"CFCFFFCFF56FC554FCFF3FDFC54DFFCF33CFEA29CCCFCFCFCFCFCFCFCCCFFFF6",
            INIT_RAM_0F => X"F667FFF4C5D45555D081C9CF33FFF9BFE5FFDBFFCFFFDA8ACCCFFF9FF3CFF3CF",
            INIT_RAM_10 => X"F000F040F080F0C0F515F555F595F5D5FA2AFA6AFAAAFAEAFF3FFF7FFFBFFFFF",
            INIT_RAM_11 => X"B000B040B080B0C0B515B555B595B5D5BA2ABA6ABAAABAEABF3FBF7FBFBFBFFF",
            INIT_RAM_12 => X"70007040708070C075157555759575D57A2A7A6A7AAA7AEA7F3F7F7F7FBF7FFF",
            INIT_RAM_13 => X"30003040308030C035153555359535D53A2A3A6A3AAA3AEA3F3F3F7F3FBF3FFF",
            INIT_RAM_14 => X"E000E040E080E0C0E515E555E595E5D5EA2AEA6AEAAAEAEAEF3FEF7FEFBFEFFF",
            INIT_RAM_15 => X"A000A040A080A0C0A515A555A595A5D5AA2AAA6AAAAAAAEAAF3FAF7FAFBFAFFF",
            INIT_RAM_16 => X"60006040608060C065156555659565D56A2A6A6A6AAA6AEA6F3F6F7F6FBF6FFF",
            INIT_RAM_17 => X"20002040208020C025152555259525D52A2A2A6A2AAA2AEA2F3F2F7F2FBF2FFF",
            INIT_RAM_18 => X"D000D040D080D0C0D515D555D595D5D5DA2ADA6ADAAADAEADF3FDF7FDFBFDFFF",
            INIT_RAM_19 => X"90009040908090C095159555959595D59A2A9A6A9AAA9AEA9F3F9F7F9FBF9FFF",
            INIT_RAM_1A => X"50005040508050C055155555559555D55A2A5A6A5AAA5AEA5F3F5F7F5FBF5FFF",
            INIT_RAM_1B => X"10001040108010C015151555159515D51A2A1A6A1AAA1AEA1F3F1F7F1FBF1FFF",
            INIT_RAM_1C => X"C000C040C080C0C0C515C555C595C5D5CA2ACA6ACAAACAEACF3FCF7FCFBFCFFF",
            INIT_RAM_1D => X"80008040808080C085158555859585D58A2A8A6A8AAA8AEA8F3F8F7F8FBF8FFF",
            INIT_RAM_1E => X"40004040408040C045154555459545D54A2A4A6A4AAA4AEA4F3F4F7F4FBF4FFF",
            INIT_RAM_1F => X"00000040008000C005150555059505D50A2A0A6A0AAA0AEA0F3F0F7F0FBF0FFF",
            INIT_RAM_20 => X"3003009000A43000026030003AAB00C0300300C330C33003300330C3030632A3",
            INIT_RAM_21 => X"C000006030030090355731832A9001900680240030002AAB30C302C3320300C3",
            INIT_RAM_22 => X"0180200000C01A000AE82BBA20022406002A326901852EEE1775001522AA0000",
            INIT_RAM_23 => X"22831809033009181A20022030C330C3158330C630330318308331833AAE3183",
            INIT_RAM_24 => X"34070000A2BFFFFC555145557FFFDB39D2E7CDCF1600E9FF196CE0BF9FE78027",
            INIT_RAM_25 => X"FFFF3C3CEAEA3FFCD001FFFFCFCFCFF366669999DF3D3FFFFF3FD407D0176002",
            INIT_RAM_26 => X"303000300A903AAB0300C0203AB20030CC3015D6333030303030303033300009",
            INIT_RAM_27 => X"0998000B3A2BAAAA2F7E3630CC0006401A00240030002575333000600C300C30",
            INIT_RAM_28 => X"CFFCFF6FFF5BCFFFFD9FCFFFC554FF3FCFFCFF3CCF3CCFFCCFFCCF3CFCF9CD5C",
            INIT_RAM_29 => X"3FFFFF9FCFFCFF6FCAA8CE7CD56FFE6FF97FDBFFCFFFD554CF3CFD3CCDFCFF3C",
            INIT_RAM_2A => X"FE7FDFFFFF3FE5FFF517D445DFFDDBF9FFD5CD96FE7AD111E88AFFEADD55FFFF",
            INIT_RAM_2B => X"DD7CE7F6FCCFF6E7E5DFFDDFCF3CCF3CEA7CCF39CFCCFCE7CF7CCE7CC551CE7C",
            INIT_RAM_2C => X"CFFCFF6FFF5BCFFFFD9FCFFFC554FF3FCFFCFF3CCF3CCFFCCFFCCF3CFCF9CD5C",
            INIT_RAM_2D => X"3FFFFF9FCFFCFF6FCAA8CE7CD56FFE6FF97FDBFFCFFFD554CF3CFD3CCDFCFF3C",
            INIT_RAM_2E => X"CFCFFFCFF56FC554FCFF3FDFC54DFFCF33CFEA29CCCFCFCFCFCFCFCFCCCFFFF6",
            INIT_RAM_2F => X"F667FFF4C5D45555D081C9CF33FFF9BFE5FFDBFFCFFFDA8ACCCFFF9FF3CFF3CF",
            INIT_RAM_30 => X"F000F040F080F0C0F515F555F595F5D5FA2AFA6AFAAAFAEAFF3FFF7FFFBFFFFF",
            INIT_RAM_31 => X"B000B040B080B0C0B515B555B595B5D5BA2ABA6ABAAABAEABF3FBF7FBFBFBFFF",
            INIT_RAM_32 => X"70007040708070C075157555759575D57A2A7A6A7AAA7AEA7F3F7F7F7FBF7FFF",
            INIT_RAM_33 => X"30003040308030C035153555359535D53A2A3A6A3AAA3AEA3F3F3F7F3FBF3FFF",
            INIT_RAM_34 => X"E000E040E080E0C0E515E555E595E5D5EA2AEA6AEAAAEAEAEF3FEF7FEFBFEFFF",
            INIT_RAM_35 => X"A000A040A080A0C0A515A555A595A5D5AA2AAA6AAAAAAAEAAF3FAF7FAFBFAFFF",
            INIT_RAM_36 => X"60006040608060C065156555659565D56A2A6A6A6AAA6AEA6F3F6F7F6FBF6FFF",
            INIT_RAM_37 => X"20002040208020C025152555259525D52A2A2A6A2AAA2AEA2F3F2F7F2FBF2FFF",
            INIT_RAM_38 => X"D000D040D080D0C0D515D555D595D5D5DA2ADA6ADAAADAEADF3FDF7FDFBFDFFF",
            INIT_RAM_39 => X"90009040908090C095159555959595D59A2A9A6A9AAA9AEA9F3F9F7F9FBF9FFF",
            INIT_RAM_3A => X"50005040508050C055155555559555D55A2A5A6A5AAA5AEA5F3F5F7F5FBF5FFF",
            INIT_RAM_3B => X"10001040108010C015151555159515D51A2A1A6A1AAA1AEA1F3F1F7F1FBF1FFF",
            INIT_RAM_3C => X"C000C040C080C0C0C515C555C595C5D5CA2ACA6ACAAACAEACF3FCF7FCFBFCFFF",
            INIT_RAM_3D => X"80008040808080C085158555859585D58A2A8A6A8AAA8AEA8F3F8F7F8FBF8FFF",
            INIT_RAM_3E => X"40004040408040C045154555459545D54A2A4A6A4AAA4AEA4F3F4F7F4FBF4FFF",
            INIT_RAM_3F => X"00000040008000C005150555059505D50A2A0A6A0AAA0AEA0F3F0F7F0FBF0FFF"
        )
        port map (
            DO => sdpb_inst_1_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_1_BLKSELA_i,
            BLKSELB => sdpb_inst_1_BLKSELB_i,
            ADA => sdpb_inst_1_ADA_i,
            DI => sdpb_inst_1_DI_i,
            ADB => sdpb_inst_1_ADB_i
        );

    sdpb_inst_2: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"1AA92BAA2AAE300024061AAA10012AEA3B03004330431AA918091A692BA431E9",
            INIT_RAM_01 => X"C00002403FFF09003003301B001A291A2EAA06AA1AAA00031A49246926A90069",
            INIT_RAM_02 => X"0018000000C0000000C0091806A40000000026003C18064C3003001500000000",
            INIT_RAM_03 => X"00190190033010010000000006E91A69001B1A431A9317551A5B306910001AB9",
            INIT_RAM_04 => X"6A2A0000F3FFFFFCFFDBE7FF7FFFFF3F3FFBC0040060FF9F1BE4CBFF35CE000E",
            INIT_RAM_05 => X"FFFF3FFCE8CA3FFCF80BFFFFCFCFCFF366669999F91B3FFFFF3FFC2FF83F3E2D",
            INIT_RAM_06 => X"1A902A902AB010002460155110002A906E90004933903ABA30301A903B900010",
            INIT_RAM_07 => X"0998000605D40000300330706EA024603AA006A02EA0181019300030AEB00690",
            INIT_RAM_08 => X"E556D455D551CFFFDBF9E555EFFED515C4FCFFBCCFBCE556E7F6E596D45BCE16",
            INIT_RAM_09 => X"3FFFFDBFC000F6FFCFFCCFE4FFE5D6E5D155F955E555FFFCE5B6DB96D956FF96",
            INIT_RAM_0A => X"FFE7FFFFFF3FFFFFFF3FF6E7F95BFFFFFFFFD9FFC3E7F9B3CFFCFFEAFFFFFFFF",
            INIT_RAM_0B => X"FFE6FE6FFCCFEFFEFFFFFFFFF916E596FFE4E5BCE56CE8AAE5A4CF96EFFFE546",
            INIT_RAM_0C => X"E556D455D551CFFFDBF9E555EFFED515C4FCFFBCCFBCE556E7F6E596D45BCE16",
            INIT_RAM_0D => X"3FFFFDBFC000F6FFCFFCCFE4FFE5D6E5D155F955E555FFFCE5B6DB96D956FF96",
            INIT_RAM_0E => X"E56FD56FD54FEFFFDB9FEAAEEFFFD56F916FFFB6CC6FC545CFCFE56FC46FFFEF",
            INIT_RAM_0F => X"F667FFF9FA2BFFFFCFFCCF8F915FDB9FC55FF95FD15FE7EFE6CFFFCF514FF96F",
            INIT_RAM_10 => X"FF0FFF1FFF2FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFFF",
            INIT_RAM_11 => X"EA0AEA1AEA2AEA3AEA4AEA5AEA6AEA7AEA8AEA9AEAAAEABAEACAEADAEAEAEAFA",
            INIT_RAM_12 => X"D505D515D525D535D545D555D565D575D585D595D5A5D5B5D5C5D5D5D5E5D5F5",
            INIT_RAM_13 => X"C000C010C020C030C040C050C060C070C080C090C0A0C0B0C0C0C0D0C0E0C0F0",
            INIT_RAM_14 => X"BF0FBF1FBF2FBF3FBF4FBF5FBF6FBF7FBF8FBF9FBFAFBFBFBFCFBFDFBFEFBFFF",
            INIT_RAM_15 => X"AA0AAA1AAA2AAA3AAA4AAA5AAA6AAA7AAA8AAA9AAAAAAABAAACAAADAAAEAAAFA",
            INIT_RAM_16 => X"950595159525953595459555956595759585959595A595B595C595D595E595F5",
            INIT_RAM_17 => X"800080108020803080408050806080708080809080A080B080C080D080E080F0",
            INIT_RAM_18 => X"7F0F7F1F7F2F7F3F7F4F7F5F7F6F7F7F7F8F7F9F7FAF7FBF7FCF7FDF7FEF7FFF",
            INIT_RAM_19 => X"6A0A6A1A6A2A6A3A6A4A6A5A6A6A6A7A6A8A6A9A6AAA6ABA6ACA6ADA6AEA6AFA",
            INIT_RAM_1A => X"550555155525553555455555556555755585559555A555B555C555D555E555F5",
            INIT_RAM_1B => X"400040104020403040404050406040704080409040A040B040C040D040E040F0",
            INIT_RAM_1C => X"3F0F3F1F3F2F3F3F3F4F3F5F3F6F3F7F3F8F3F9F3FAF3FBF3FCF3FDF3FEF3FFF",
            INIT_RAM_1D => X"2A0A2A1A2A2A2A3A2A4A2A5A2A6A2A7A2A8A2A9A2AAA2ABA2ACA2ADA2AEA2AFA",
            INIT_RAM_1E => X"150515151525153515451555156515751585159515A515B515C515D515E515F5",
            INIT_RAM_1F => X"000000100020003000400050006000700080009000A000B000C000D000E000F0",
            INIT_RAM_20 => X"1AA92BAA2AAE300024061AAA10012AEA3B03004330431AA918091A692BA431E9",
            INIT_RAM_21 => X"C00002403FFF09003003301B001A291A2EAA06AA1AAA00031A49246926A90069",
            INIT_RAM_22 => X"0018000000C0000000C0091806A40000000026003C18064C1775001500000000",
            INIT_RAM_23 => X"00190190033010010000000006E91A69001B1A431A9317551A5B306910001AB9",
            INIT_RAM_24 => X"6A2A0000F3FFFFFCFFDBE7FF7FFFFF3F3FFBC0040060FF9F1BE4CBFF35CE000E",
            INIT_RAM_25 => X"FFFF3FFCE8CA3FFCF80BFFFFCFCFCFF366669999F91B3FFFFF3FFC2FF83F3E2D",
            INIT_RAM_26 => X"1A902A902AB010002460155110002A906E90004933903ABA30301A903B900010",
            INIT_RAM_27 => X"0998000605D40000300330706EA024603AA006A02EA0181019300030AEB00690",
            INIT_RAM_28 => X"E556D455D551CFFFDBF9E555EFFED515C4FCFFBCCFBCE556E7F6E596D45BCE16",
            INIT_RAM_29 => X"3FFFFDBFC000F6FFCFFCCFE4FFE5D6E5D155F955E555FFFCE5B6DB96D956FF96",
            INIT_RAM_2A => X"FFE7FFFFFF3FFFFFFF3FF6E7F95BFFFFFFFFD9FFC3E7F9B3E88AFFEAFFFFFFFF",
            INIT_RAM_2B => X"FFE6FE6FFCCFEFFEFFFFFFFFF916E596FFE4E5BCE56CE8AAE5A4CF96EFFFE546",
            INIT_RAM_2C => X"E556D455D551CFFFDBF9E555EFFED515C4FCFFBCCFBCE556E7F6E596D45BCE16",
            INIT_RAM_2D => X"3FFFFDBFC000F6FFCFFCCFE4FFE5D6E5D155F955E555FFFCE5B6DB96D956FF96",
            INIT_RAM_2E => X"E56FD56FD54FEFFFDB9FEAAEEFFFD56F916FFFB6CC6FC545CFCFE56FC46FFFEF",
            INIT_RAM_2F => X"F667FFF9FA2BFFFFCFFCCF8F915FDB9FC55FF95FD15FE7EFE6CFFFCF514FF96F",
            INIT_RAM_30 => X"FF0FFF1FFF2FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFFF",
            INIT_RAM_31 => X"EA0AEA1AEA2AEA3AEA4AEA5AEA6AEA7AEA8AEA9AEAAAEABAEACAEADAEAEAEAFA",
            INIT_RAM_32 => X"D505D515D525D535D545D555D565D575D585D595D5A5D5B5D5C5D5D5D5E5D5F5",
            INIT_RAM_33 => X"C000C010C020C030C040C050C060C070C080C090C0A0C0B0C0C0C0D0C0E0C0F0",
            INIT_RAM_34 => X"BF0FBF1FBF2FBF3FBF4FBF5FBF6FBF7FBF8FBF9FBFAFBFBFBFCFBFDFBFEFBFFF",
            INIT_RAM_35 => X"AA0AAA1AAA2AAA3AAA4AAA5AAA6AAA7AAA8AAA9AAAAAAABAAACAAADAAAEAAAFA",
            INIT_RAM_36 => X"950595159525953595459555956595759585959595A595B595C595D595E595F5",
            INIT_RAM_37 => X"800080108020803080408050806080708080809080A080B080C080D080E080F0",
            INIT_RAM_38 => X"7F0F7F1F7F2F7F3F7F4F7F5F7F6F7F7F7F8F7F9F7FAF7FBF7FCF7FDF7FEF7FFF",
            INIT_RAM_39 => X"6A0A6A1A6A2A6A3A6A4A6A5A6A6A6A7A6A8A6A9A6AAA6ABA6ACA6ADA6AEA6AFA",
            INIT_RAM_3A => X"550555155525553555455555556555755585559555A555B555C555D555E555F5",
            INIT_RAM_3B => X"400040104020403040404050406040704080409040A040B040C040D040E040F0",
            INIT_RAM_3C => X"3F0F3F1F3F2F3F3F3F4F3F5F3F6F3F7F3F8F3F9F3FAF3FBF3FCF3FDF3FEF3FFF",
            INIT_RAM_3D => X"2A0A2A1A2A2A2A3A2A4A2A5A2A6A2A7A2A8A2A9A2AAA2ABA2ACA2ADA2AEA2AFA",
            INIT_RAM_3E => X"150515151525153515451555156515751585159515A515B515C515D515E515F5",
            INIT_RAM_3F => X"000000100020003000400050006000700080009000A000B000C000D000E000F0"
        )
        port map (
            DO => sdpb_inst_2_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_2_BLKSELA_i,
            BLKSELB => sdpb_inst_2_BLKSELB_i,
            ADA => sdpb_inst_2_ADA_i,
            DI => sdpb_inst_2_DI_i,
            ADB => sdpb_inst_2_ADB_i
        );

    sdpb_inst_3: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"4000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000001004000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"BFBFFFFFFAAAFFFEFFBFFEFFFFFFFFBFBFFFFEEAAAAEFFFBBFFEBFFFEFBFEFBF",
            INIT_RAM_05 => X"FFFFAAAAFEEFBFFEFFBFAAAAEABFEFEFEEEEBBBBFFBFBFFFFFBFAEFAAFBABFFE",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_09 => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFBFFFFFFFFFFFF",
            INIT_RAM_0B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0D => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_10 => X"FF0FFF4FFF8FFFCFFF1FFF5FFF9FFFDFFF2FFF6FFFAFFFEFFF3FFF7FFFBFFFFF",
            INIT_RAM_11 => X"BF0FBF4FBF8FBFCFBF1FBF5FBF9FBFDFBF2FBF6FBFAFBFEFBF3FBF7FBFBFBFFF",
            INIT_RAM_12 => X"7F0F7F4F7F8F7FCF7F1F7F5F7F9F7FDF7F2F7F6F7FAF7FEF7F3F7F7F7FBF7FFF",
            INIT_RAM_13 => X"3F0F3F4F3F8F3FCF3F1F3F5F3F9F3FDF3F2F3F6F3FAF3FEF3F3F3F7F3FBF3FFF",
            INIT_RAM_14 => X"EA0AEA4AEA8AEACAEA1AEA5AEA9AEADAEA2AEA6AEAAAEAEAEA3AEA7AEABAEAFA",
            INIT_RAM_15 => X"AA0AAA4AAA8AAACAAA1AAA5AAA9AAADAAA2AAA6AAAAAAAEAAA3AAA7AAABAAAFA",
            INIT_RAM_16 => X"6A0A6A4A6A8A6ACA6A1A6A5A6A9A6ADA6A2A6A6A6AAA6AEA6A3A6A7A6ABA6AFA",
            INIT_RAM_17 => X"2A0A2A4A2A8A2ACA2A1A2A5A2A9A2ADA2A2A2A6A2AAA2AEA2A3A2A7A2ABA2AFA",
            INIT_RAM_18 => X"DF0FDF4FDF8FDFCFDF1FDF5FDF9FDFDFDF2FDF6FDFAFDFEFDF3FDF7FDFBFDFFF",
            INIT_RAM_19 => X"9F0F9F4F9F8F9FCF9F1F9F5F9F9F9FDF9F2F9F6F9FAF9FEF9F3F9F7F9FBF9FFF",
            INIT_RAM_1A => X"5F0F5F4F5F8F5FCF5F1F5F5F5F9F5FDF5F2F5F6F5FAF5FEF5F3F5F7F5FBF5FFF",
            INIT_RAM_1B => X"1F0F1F4F1F8F1FCF1F1F1F5F1F9F1FDF1F2F1F6F1FAF1FEF1F3F1F7F1FBF1FFF",
            INIT_RAM_1C => X"CA0ACA4ACA8ACACACA1ACA5ACA9ACADACA2ACA6ACAAACAEACA3ACA7ACABACAFA",
            INIT_RAM_1D => X"8A0A8A4A8A8A8ACA8A1A8A5A8A9A8ADA8A2A8A6A8AAA8AEA8A3A8A7A8ABA8AFA",
            INIT_RAM_1E => X"4A0A4A4A4A8A4ACA4A1A4A5A4A9A4ADA4A2A4A6A4AAA4AEA4A3A4A7A4ABA4AFA",
            INIT_RAM_1F => X"0A0A0A4A0A8A0ACA0A1A0A5A0A9A0ADA0A2A0A6A0AAA0AEA0A3A0A7A0ABA0AFA",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"4000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"BFBFFFFFFAAAFFFEFFBFFEFFFFFFFFBFBFFFFEEAAAAEFFFBBFFEBFFFEFBFEFBF",
            INIT_RAM_25 => X"FFFFAAAAFEEFBFFEFFBFAAAAEABFEFEFEEEEBBBBFFBFBFFFFFBFAEFAAFBABFFE",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_29 => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_2B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_2C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_2D => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_2F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_30 => X"FF0FFF4FFF8FFFCFFF1FFF5FFF9FFFDFFF2FFF6FFFAFFFEFFF3FFF7FFFBFFFFF",
            INIT_RAM_31 => X"BF0FBF4FBF8FBFCFBF1FBF5FBF9FBFDFBF2FBF6FBFAFBFEFBF3FBF7FBFBFBFFF",
            INIT_RAM_32 => X"7F0F7F4F7F8F7FCF7F1F7F5F7F9F7FDF7F2F7F6F7FAF7FEF7F3F7F7F7FBF7FFF",
            INIT_RAM_33 => X"3F0F3F4F3F8F3FCF3F1F3F5F3F9F3FDF3F2F3F6F3FAF3FEF3F3F3F7F3FBF3FFF",
            INIT_RAM_34 => X"EA0AEA4AEA8AEACAEA1AEA5AEA9AEADAEA2AEA6AEAAAEAEAEA3AEA7AEABAEAFA",
            INIT_RAM_35 => X"AA0AAA4AAA8AAACAAA1AAA5AAA9AAADAAA2AAA6AAAAAAAEAAA3AAA7AAABAAAFA",
            INIT_RAM_36 => X"6A0A6A4A6A8A6ACA6A1A6A5A6A9A6ADA6A2A6A6A6AAA6AEA6A3A6A7A6ABA6AFA",
            INIT_RAM_37 => X"2A0A2A4A2A8A2ACA2A1A2A5A2A9A2ADA2A2A2A6A2AAA2AEA2A3A2A7A2ABA2AFA",
            INIT_RAM_38 => X"DF0FDF4FDF8FDFCFDF1FDF5FDF9FDFDFDF2FDF6FDFAFDFEFDF3FDF7FDFBFDFFF",
            INIT_RAM_39 => X"9F0F9F4F9F8F9FCF9F1F9F5F9F9F9FDF9F2F9F6F9FAF9FEF9F3F9F7F9FBF9FFF",
            INIT_RAM_3A => X"5F0F5F4F5F8F5FCF5F1F5F5F5F9F5FDF5F2F5F6F5FAF5FEF5F3F5F7F5FBF5FFF",
            INIT_RAM_3B => X"1F0F1F4F1F8F1FCF1F1F1F5F1F9F1FDF1F2F1F6F1FAF1FEF1F3F1F7F1FBF1FFF",
            INIT_RAM_3C => X"CA0ACA4ACA8ACACACA1ACA5ACA9ACADACA2ACA6ACAAACAEACA3ACA7ACABACAFA",
            INIT_RAM_3D => X"8A0A8A4A8A8A8ACA8A1A8A5A8A9A8ADA8A2A8A6A8AAA8AEA8A3A8A7A8ABA8AFA",
            INIT_RAM_3E => X"4A0A4A4A4A8A4ACA4A1A4A5A4A9A4ADA4A2A4A6A4AAA4AEA4A3A4A7A4ABA4AFA",
            INIT_RAM_3F => X"0A0A0A4A0A8A0ACA0A1A0A5A0A9A0ADA0A2A0A6A0AAA0AEA0A3A0A7A0ABA0AFA"
        )
        port map (
            DO => sdpb_inst_3_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_3_BLKSELA_i,
            BLKSELB => sdpb_inst_3_BLKSELB_i,
            ADA => sdpb_inst_3_ADA_i,
            DI => sdpb_inst_3_DI_i,
            ADB => sdpb_inst_3_ADB_i
        );

end Behavioral; --Gowin_SDPB_8k
